PK   y�:Xp:�  ��     cirkitFile.json�]ݓ�6��W��������ݫ�î]���R�$�"KsM�l����'	BjMc<q֓�x�hv7�n4 ��dcq�y�޸�/n�X�&wDL'��dϯ����b5߮�?m��������b�۽+�����ʭ��TH��ئ�Tԅ.�-���U#X%H;/'wo�O�|;��Nq�3����>vsk[���
�,+xMTaJR̱��e���'GH�%F�LH�sF�M!]���Vڰ�h(�J	]kJpϬ0��0�uB��:�Ia[Zܕ�0̚����+�hŸ�(B�AzW�мT�ReD��)8����g�X�W��[��	!��B�PFq�YB��������Z]pFL�5��-�4�q��Ft*�D��:�@�qO�#�hTT ���
�$�@�J42$Qd�@�2e�Ȝ��ܴ4ι�i��H?��)*Y��:Q��Y��8�Д��D�|���4�:妠�)*q�=5�M�M�M6�G�
cz��p�h�P��:CMp�U+��'a4`څ�J��	Bt*I�f|�)߄f|����6���
�� D�FPh$N�6,&aD'3]X$ƈN�`��MQ�Q�ISN�1O�K��B4�Q]��i`I!95� G{�g��?�����Cw2-��0���l�	')��n�)��nѩ4XnF���?����r�A.M�Zv?�
Q.4���qi[�\D��l[��"-�A=�
\|f�Cpс�qe�1Od�n^R�Ra�t�U�6Ű��۶�q�a�vlS�=���æC��c�u�a#wڨ�6�Ek���ޙ�����Ƀb�'�L18O�y�0�P�:�}�C��Pa\�v(vZ�
?ڡ�t��(m�(v�Ą-��,�Y�L�D�b�Y�0яu(�J(��f������C,�Y	���fbh]��0-�^����c�pzy���@3XW\�U��	�@yŗ���+> ,^qH`���,�]��u��9,��vy�-�]�;AK_��+�2��`�H]��A�KW&�BѕI��s9���o.g2�J��DZT9�LO����:l�d���DH�\h.,�����Efᢲp�Y��<���<�%y�K����0Ƀ`��$�I�<(�yPL3��<(�yPL��A1̓b��4�i�<(fyP�2�yP���A1˃bv��	��UԀ$x.W1.��\E�@��r=�A$x.���@��r/�	��U�$x.W�.��\}"p��2^�<��O.�����ܺ����_���#�E���O'��0�_��5��j��4n3�{��5�0Ĳ��B��y��M�mE��J�h�$�ۿ��N�t�':��]�D'@�N�D��8щR(H4y��_&�3�ˤ�a~�4?��/���e��<����>5Rtb���0�E���k��}-���ڝ}�M1�q����10Í\���	nGFtb� ���U>��6/f�d�Z_��o��&��CC��6�ۢ��rB2��Z2�<tbF>�.}|
�N4���Z�ǈF���cvua$��]I����������q��k�vՌ���Jz��ߗ[.�4xA�Yl�\�Ƞr�"��U� 32h�\����{_xA�5�v^,�`��s�D�"���D�Z���D����D�����D��3���,����%ɗ�A�<��� �r��v�6����H�q@mσ�,6�i�\�E���b��9l�� ����T�'W/d�N�3�0l�\�2� � ��� Wѐi"V:�~��,yj|�R��gS �a�y\�y�),�r��/;�yB�7|��7�A����(����
 w�]T��l>Û �����@��=�������s��|��qx�;�.j�%6�����k��66��M�X� <��>�E(|\4��	�� �����pL��I�� ��;L!S���0Q���|uȎb<�`�XƏ��t�����@c~��N���s�/��獝u�<����8�ݡD}�"����
�CPlp�������1A��DxT�1�1�������?��"P>�j��YF7fXg#G}�a$pc*6�qL`�NFLt �L���%||8�f�o�&��M�q�v�_i�la6&���^��)τ�t$詊v��X��654B�Y�sK����0���A��G0�a��#�Ô�F6�d���0���A���R0��8`�p2�	�}v�||����ve8���fф*����L��9|�48~x̠[p���6���EC'u����Kv���CY����n�J�	���n�`�W��;h���;h���;X��u�;���ݞ[�`ݗ`!#���� �����u_P�Ċpc��<��w}Ճ4������o(/tk\��p��e�x��8'����x�=���rۀ��^����c�a�qڈ�{�b�&b���g�m��4�9F�a~qʋ�{�_��b�Վ=�/ΐ1�`��l�6�#�����q��uqz��{�[<;�����8}Gh�=�(�� ��fϓ�`�7��E��|�#��Y�4�S��9Ɵ���s��6_���x���}�Q<e��k�nʠO:�'�m��8NS�m�X��Vn�͢?~�O��Kx�A�7����h���M,n��&7�}����I�Mjߤ�&�o�q��7����Abs��9b{��=Hlr0�-B!�I��$$�	9؄�F!���*�`���Bb�Ѓ]hlz���B�8���c��y�q���v��j����a܄��fֶ��)�hJ�	���T*Yg�\����7�����K�n��%X�?�$=��n���{w��f}�6ۅ��J�W��g^ۇ�f���?��~�����|�W�X�x���2�=|Xz����ܵv��|����xXTKw��q���ظfr����Ѯ[[o7����dg���ce�$|ov���.��o	Q3?��R��PL	3I���Ľi��?x��6�Z&Q����ｦ��p��]��L�1�X=l�����M'������i6y����Ŧ^�}o����L��M�)�O�RNg\�u� ԌSCN�1�����fLH�����������جT��k SB��J��:�@F��d��8AscfƘ��@�ƹ������ƹ���<����������42�	=���#�N�q�Ϙ�vI:��e�s2�8��Y�q:�g��{��8�f3ͼ0q�Lzn�Խ��8�`3C�������p��򣎠q�n��t'?o?9�x�����c�#t&��+f"��SA�+�(}ӄe���:�����L(���ԇ[�O���c��d��3��؞?4H5��I��7����w�*4���ϋ��c�X��6�XHfd�ԑ��Ai��P�pfZx�3-<��N=獰��sRh�d�����O*|�&֧�ƻ��s���0�w��0���t��A]ozo���n赐S��ƎMe�SS9+Ǜ���N>;oxG�J(� ����ʙ*}>r�rVΈ��8���>gN4e�:?��Ͻ�����7�peńk%��p�2`�Q�p<b�:O\��oa,*�	"��`O#�˘&��n�V���~bW[���εE��O��K]���Ȑ�e7�!��b�u0���!��I<�i�h�$ޔV�ϫ�
B����ͽ���ߏ�왵�hԂ�r�^��[>ݖ'��Ebn$�\��U--���5���+J�V��D�&�R, L2��T�~tR!��Z�8��D�ip���u��_�SW��(���zi7��og,���LϮ칆y�Ŏ��N������D�����b���Qvw�צ���?m֏������3�N�iNO�׶������_�ۺ��cBTG1�"�PFJ�~j=�z��Z�������n���Ȕ^V2ܐ�t����G�����}��^߃����'�Z��+���Dť"FNz3�2J
̘�!�C�f�$��>��s�hf�q݁�c�a�r���!��D�����umd!��hUT�&�TV�u��*J �: �*$�^A��r�}~>ކ7�sDS2�ͳ�U~�7��@�V7�aE#y�,,�n*�Kɪ�WC�6�@r+�3 �ң�z�-���+�>��-�(�]�88)�
�r�e�]��	��g�&�/���C`A���RuO?��O��U�g~<����[_@�f����X�{�q��o?.ܧ���C���w��k��&w�B�4L�w��;?�؍ʫ����{w:nn�\���ӱ��Oo����=�z�����C���w��MBY�U�:4���p��m���3?�����MAzS�#�`Ju?Ow����&�=����uγ���CG�<+:�'��W�K��O���3w���ӁdPl��,�*+6D>l���Y�A���^�7��>M!�N��$���T"+6d>l��ؐY�����^Y?��>M��:�7��ɠ��mxތC��ɍ��)��-�$��+��h
����H�Oۖ�4Y���G䆏�
�����ơ�')��h�_* �A�!5kXք�e�ʨ��`y�2�I�No�oNͨ���E(<]��:Eh:���7�� ��w#:z�LsN���[�R�@�s���e�>���g�s���y�>����T�>o��7��s���i�>'Y����s2Z�bO�*�:�ù�j����G	�+�=��&Nf�S�[�ág�/YoHU�Q��vi�@D��MC��M`���S�	8�ܠލ��oʜ�wd;���X0*>>=�v~\���wEfXNh���W�2#\�A;$0zۈO]�/B���xAl��jNȶ�Z�U�a�f��~�v���)85gP11J�e0*>^k�'�JU��V����77��'w1�>w�v7§�W<���]��+o0��v�$|"��B�?Ykf���{��kf���Ի�f��מ�������WJaTzT��M�b�q�hao�l�^�·���'/x�}��*��!U91d��Q�DD���8x�{�=z�ϖ��Ի5���MK���i
5:=�F5��%�f-\N�Agd,�ܲo�[�B����%˶�u]6�!߅��V��^)UNld\�!�$5p�ra�<-�,槰1\�OO�n'KTu��aD�X.te��N�a�`G�d���n����^�>u���k@Ta���Ċ����d���xm��-V˃�̒\̻A�['ݴ_g�[4a'�h�v4�d�dՉ2ki�f��:4oDxZ����{���4�76 ���:=���X._���[�Y����.���c�o��î�������CP������PK   �{&X��N���  L�  /   images/3e5d0cfe-dbb3-4add-86f8-df5e0b35ef62.pngD�cxf]�-�IǶm;�ض�ƶm�N:�m�N:�m�����s��Zk���ԬcԬ./+����/X	qa�_��/~�� �~�J���?/ GE1�_��8�?GA	e��0
���������[�E�j"����3�Tu�c����*�iȀ���*R��|�]�Iϩ ��ڇ�
=T�m�DB
�|������V���u���魐*j�?ج��/,~T���qǻ����׬�kנ�-G��gu�6�oށݸ������x�����&5����e��r���g7FX}[�we>W���[��-�T�a��Sy�¬��f��)�D���=Z��s��cW��g�Zn�������^$�½�x��h痎�y���8]�#�]�*nl}W�\j�**	ƘKk����k�c����Q�@`����a����u1חĚ� ��{���&|Ү���?8*�`C~l����6f쿉��q�on{o��<���r*�nJi���dV X��(��.��VF�F1�[�K�xd:�]�K�e�=v�Ӏ��x�^�F'wkç�u�t�(������l��l����|���ԥۍ.H3����!���~g�YwlS �N�-K��xH�X��G;ĳM=6/�\�e�@!lX?�4�[��t�(��.�?>��~����  H[~^]Vі�|Z��{����Kf����Ѯsԏ8���g6���ҷG�]Ty{`sh~?�6�ٯ]�I$�������QN���u��֮�9Z�w�f*�0���N��o�D1��rVn�w��IO��[��yWG�{4K�9��;,c��e����~��x�K��[yMë �S~���2E��g�ex>K�饞�-�(p,���Д2� �����5�q5ۚ3�h���2��HEx�̳��)�Д�B�TAf��b�F�;?���]nԱ5=:2[�3�1���;2K��� �}Ƀ1��t����<*��E���|�)e���V��`��EK'���|���ߧ;���Ţ9�ıHH,�0C��,�騧J�-Ii�>*Y:��� |H9���8�X�HY^��^��bו���n�9k�\z���F���3G���{�T8�X?y�6�8�cU���lh�R�}����IU�ߊx�
�ܾܺ�5����3����5��X�qi�������B���@uv�T�ֳu�T<��+�u�ʉ�č#�a�?-��NK�D�M�g5��2�V�4�Z���a(K��^Y;�	��)��s��p�m���u�Gy��}/^:�L���%!����C�,�-gY<���ϷEW҄��|��$��I8�H��p��a��p�F���G����Kֆ�gu1���[;Irq7�~[U&�v\ڵ��S��(\�D
�O�1%"�����3;p����*��;�����Y+A��Z�Y+	p�y�h��Ϯ��5�.[7���f�mD�T�VZ;�>>��v:�:����G�ٽ��u�����>]��$��8K-��9��s���X��j��{��!�ך�k0����nl������:23���}���U��;�}�#[Q���Μz��..���*৊���D�X\��^�4���.�ql�{��|U�I7���B��4oV5�|����$l�7�q\Z~��zu{7�&:1��z�P`8�6����I���m_����d�Bg*8�\c��A�Ƃ�Ɠ]'������
d�p�|�:�>�q��x}\7�:��N����WrW��H�!��2��5W�	~��m��p�u@�M5I��lEc�����@O� �M������:�P���e�0����$�qhޔ�*h���1�m�� �!�wwb�����]͂t��[Jɋ��=���8#���V��k9� �~t��:o���:/�=��4�[�5Ra9�ֻl���v�Z�{���T|&���'f@�a��/)����n#Ln���ιgnBBP ��������CT����쁷�[G��A��#M�������̖D�����g�kjkNo�W��R�v$D��DH̴�����k�����S�H(��y��,W�^/%b�hTiBݳ���tޜ�����CG��q�8q&K(('�Q@�s(Ǿ���������U6)�q|�t�c�l9�y	�BD̃GT�*��џH��1¬��uv��L�#c�����$�ݲ�;g�t�yd-���G���� �u7 �s�.'�L�-�}X9$b����%e��xn畬I�ys���*�8qKv�L^O\�H�0��)2��uݏ��dc��m�Q��
B�LC�4,��k�ڻ�����VQ��^�x
iI�q�:�G�T������F���F�ߺTP��s�3�N�>��v�ABW�V�p��:��@!V��2.�QQY�c.1�n3C��>�����	�[�u�I�mv�z�p�K�PR`��D �Q63&�<�O�o��|���z�0�ҕ�=��ln�fLSL@-����-���  ��/��9V0�5�@D��b�����VS3��բ:��=a���6G��{��:��c���v�W��?E��h\�����LOW���v��0����c�6N2��5b��9��b��<�z �8ł���/�t�ш�)E0�țP�$�LE;e�D13�Gw^�K�30����L��*!�3�����qOXP:�3t�$�n���Qh��s�t�n��w����Md�<7n�z�q�(Ps�����{��q&���]6dm�ރ�eo�����k��.8_�qW���{�f�^K����J�}&Yqe�E��C���\m�]��_�~t�/4�V�����c��: �������'���}ε����.��_i}
�3��h@ �Eh�T��c�{�8���d���w�u}=� Յ˭��s3!a�w��Β��)67_�����$Y_S��C��e%)g��.�<R�C$7�(X�ҹ��WL0̸��h]�fِ)�F�������Y%��%f~�j{i�Pz��v��j��M@#)�]b^�n)afzL6�V��\8=k����xf01i]S�:��^�*iJٱ��i���yF�oNd+��v��S����ChQ�,� � \Ң��\���ݣ��h��[���ʭ$:OExi�n� �߈֏��F'Z��C�Y��L�L`@v�Hҝ`'�`C9n�����i� ahV���۶�i�����Oq��.'�� ����u ���Q�7�E$D�,y�WqŔ�8=���
1E��5�"���}5�LS)�H]t4_�8k%�9�ى���j*i4ĵ)zِ��P�0� a"�u@$#�a9��SB�\}-���*��"9�4G��o?��"�sSN%S�VlZ_��ﾆj��/D|���C+jm�j:ޮ~\+�?+�.��%���Nq/��_��4��Dy�L�!���R��N�q�����/�t���~w��Ơv���Lo���^��*$���]�qZ ᑹ��7�����.TDgn#sO��y�����VT0}r9s4�'��+��x���/��O�D�~C��5&�ϟ�Y4��nբ�\�d�V��a��7cNL/��5�A�
�����S7�����h�9e���VM�l��18�8�%/�@��&�j�-z��0�/��5�\Zϟ�J�&���)��W��Xсwv^��[�ˢ4�Ɋ��yh$�<�֐h���LH�����Q��c����s���ͭ^����I�ԜĦ[�d\9�*õ������Fp���1i<s��87i]Vo�<K���A��iEHmBص�F��9<����tUȂ�۴A��3���\o60-3Ob̍�8�����V�;T�~BA'pLMr`�Â	��z8�3�Eg��7�����`"L�	s3d�q�SOfmY�V��=�TO��tV�C��#���� ����n�S��T�]&�v��]�]H����	��#���KF�_��<"<�Fڈ%�6[\�#�򼃶�l��f����E(��H���L���$}9~��ۣr-x�V�q�?V>	p�Pߌ3G�_(Ç�"
B"ýy�y��o�	��O9Y;�-�O���4�HƘ�
��L05R����l��9�����vS���˩�U:*JWQ8�����➸�s�N��%h�n\#�^���R��y;y�}X��妢�B ��ٹ}�OV��-o+r�:ט�H�q�������X��R��J���JQ	q��w�L?ʾ���/�W()P��N�������¿��H�D�DH���{h^gh��I���J����`Ы�gW��|T[�
����g�3��nQ~��`���U�r\e#sӠ�}�b�` Ҫ�V�7=��r���,�P/�Y�����3�_�u�r��^h�v��ʝ,B�Y�*)Ūl�l��bZ� �2GJ>.t�y�SR�1̿3��5%y�N�hd�B��&XY��{�L\Uc�[*"�o�@��@�8,Mb�U�'������~^W�OA�/5�P��@KuI/�a�d���1zy��3���{����o?u5��ơ��NEOjV���UL��Y���	s�F�� 7�h�躢\q�!��z�p���h�*�Hp�PMUj�/4�>�c�;�����@����ZEQ�p��YR��ݧ�K��0� '�fR��pGF�o�����C��I�:q:qf�!���G��bē����u���
�.١��a&͙�g�p�V��#�Hx��u�-�%b���
�8xT��|�{���[��v�XR�t�?E��؎��<�'��;PeY1K6#���p�ψ�[/M�B�?+�ب1`��|U��~HD7:Xxw�������J%ѥc��}�]��>E�G�cKL�|�������"�fD����lT���L��yyl�14S7��A��RGN�_�����s���Kl@������WD |ѥ��!¦'���#Q�@�`���ɣ
��(���u�dɘ�=2�����d���C<L��K���U�;�P�ޭ+{dbZIsIn}�w���l(j�[�`�p�t���ӹ�c-h)�D���"�G1f�`���T����y��{�!`,_,�)4�5V����? ���03ۀi�.E>:�����{a���c�� ����
$���C�Y�tEx�a'��x��r!���Kl�/�T��;յV��Љv���@w�*+�pQ$��ٚ����G<�N?���G��1<�c^���p�B2y�>���ʣTb��Ǿ�ƭ6��������.<�
����iK1�ٞȴ%裃Ϛ�C5>b@�/��݁�x�Y�z�a^CW~�	NЙ�n	����rZ�ٌʠ��.�~���*$2�(�۰��j��n|��(�e�֙�Kl\V�*��T
v�;�}t����r¢zR�\� ^B+Fx�����n��P����a���M}jj���^��Z��3�b&I�l�'=D���ڍ?ðG�yMś6�J�)�I�Y�Q����V�{�(p��n��8�1b�}_xg;���;}�7������N^(����v��$?֠l�A.�K(E*�������� ��9,�C��Q@�k��(L�����u����}�lR�`��Q*A���G�K爌�5�=\��_�1�a�Zy��Oj�=�V4�6����֨.]�狝�0l!�w�`�����9Z�8������Є���7J^�4_lz����fb��,����W���d����B�r�<����Y"!Ju�\�ٍ��C�Zڪk�R����ZGG��U��`|Fa�xK�&OE�Ъ���c]�<Ah�}W�P���$� �� <�ꠌN�G�uWWv|�p�C����WY�W��ib������x���S:�Pb��r���ۀ����1��kS�;cW��|7��>�X�gW���7��3d��[#�QR�Tw��D�eS�@��F����3�
I�a�rI_KǠyL��^0��$�̜B�������?``�!��Ɋ9yTM��N}\�F��v�50��I'�qH� �1�r���c��4�
��l�o�H�������זTT;�"�+�E��`����ei����y�o
�s����ⷴwG���� \�S��&�0W���Ez%S�_:��' �~+�y�"#S:��\�_�V�bG���c,���6�S��}�[�O4.-Vhq�>�1L��V��lImV��BzT��-@Ro�]�����n4<gwT����ӹ$N)���x��p�U�� "�_�^@#Y^n`bjdՄv�����h�9$gJ�uvv��G�)J�p�g�"���-�re����S&C�ְ�DV�~��"�5�@�kT>���CŔt�Ƀ �3k��%!��h�G9]='uI���,�a�XC �Etܧ�,WF�5����&+
��_"VU���;�ĐߒxbV#�ݠ�����Rq���(��)1��{�������+,�g����TP�Fz4�Tt�5�^Bf�wa��1�����s�"UV��DMEЈ8�Ao�w��ҸQ4�����-H�_���|O(to�6B�VjЖ�M�/��rSL$�R�����H������۳�ǌ���8���Z�Ex�������8[s�x$���L��Q��.��tm'Y�N���WBQ/��;	Y��̙R��������-#՘�'|�oBdn�
�pMٙO��������rO|J�P�Ƴ��w��g�MP�� Jg@�Q�R���p�RR��"�%�ٹ�n�Ԥ/k�}�^�ވU�����$p�ԏ��SNH�x[G�șS;��
��&�=�ԅKYeȉ���&�5ᗂ���6y�o��;/�` ��&�=N�������Ǔv�#:-vP�������m0��]uX2��mJ*I+I�0$YD�b<)�1� A�w�q�Pqj$��sn�.�~]�fP?:E��)
%� Կ��4پ�QmY�ä�A���'������'n��Cv�ՉwqB�6aB��E���n�A�3G�3u����~��}��7���O�qf���g��t��Xk�\�������3�ӥr2�~ī��%T���c�����-�eI�rh�#��dQm���t^���J�P��|�ѓu����\<"�����1�{��'k <�V����N�0�r����͵��5"]c���h�AI�"�g�ǭ�袻l(Iֻ�<}�BUFS���	g̝}�Ҕ&����H��2B�|t�Ո�0C�� ���I7!��%M6C��CϜ���r�p)��
'��q���[��-f�Dcއ9x �25�.�~8�*�����B��LOd��V��1]�o�+���Zb�B~�,2�M��7RK��u�/_-��n;����'"�-����F�W�yݯ��#�Z4}��gnjI(��^+�~��K��ʸ���5�5����$ll�K6���z�p+����~�[��m/X�Tt���Ǚ�$\�æO���-����BK�U�d�|����ll9�=S#�5�I�o̟��bcSY��ܒ�=�����F�cl6���P��>�.{v���aӕM�o Y�v���eJ%�#ul�|�0U`~䖗#I�Wѩ���yz��Ízy�&%>0�s
�������lS�l�ߤk^p�Lc)�@.^�곶A�rk�w��&w�"���d���A����Z��x	1m��,�׆�Y[T��g�0� Fc\?:j�q�myݫjC����>�6��m�?b2,�HLS5+9�pO󿩷����C79���x4�x�;�'1�?Y�Xg�|��&\p�Hy?V�p'��Od-CU���,����"��F��QD��A�V{�h���~@9ߣ9xfl����n����Y
�^�7�k��/����0�Nw���t;D��EW/��Ŗ糗H-Jw��gR=�mg�XtX��p���8	�H��N*�)���A��ˆW�wT|���Dz�_��>���e��Cy<��P�J1�!��ɟ15��7i2� �g����*��\��>.PԐ��$9v=��A$Dy�n�3d S��~p�������b��X��t�����S�>k���i�qя�*��mߧk!�!a�,	�����L$	��^	����Ս��'�A�r�|��E1sɨ�_���uU�	A�ɨk���]�J���.�h�-�H�a��:�É��E��Aߏ�����x�?�3�K�])��/c)�u�u����Ϩn��~\��)hi�Q�G���¢GB��Z�������/HQ)�w���U�t-^���Qsm��Dו��|��~��-�*q�?e7��H(;�_C��0�Ine_�% V���\E�Η����R�_�H��eS��gT�F���A$(:��.� ��8��<az�q^U��d���;Uu����������i@H3����}�vh�9;$=�0�KeU��+z���JٵM�g<.���gJrr�p��W���j�$����p��  �s5n�i�ģ�B��K�z���1�S͐��ܵpw���\��-�
�1a�M��.�շ9$Fx��<M�biy��WYE��Cw����%��?�R�*H�Q�w<\P���W�������ho�ζ���nJ��S/���J�S@'Mi1��@{T4|�E�0q�s�9�P_f��1Y�YB��4�r�:�C�x��k��+�Oֆ��_�J{��e�4E�����h���vA��M��?�"��óp�i�l`��!���8+@LCԅc`�s<K�p�1i(�WҶ�\�!n���T��(Z9�q9��$V.K��9>�mR���[� ��"�H�@��<�3���4xuَ�	�`'��B�\�8؁9m�5޾r����]�^u��]�~�����O�<U��oSߜLk����b��� �h��X��#��W"�!cj�����=����mX�7��<BFI\icj�������H��Yc�ߙ�*Hc�?n'��uC��@��mU����Ƽ#K'C�s��D��	sc����Ҍ���}�F�che3;�(S�hu��d����3���Q��D�7����S)^�l� zm�SI�(~:V�W������v(�$RT��Z�n�����d�U�E�`�>%v�>��Wά�@8d2�9)�A�S��]2��
���V� �$M�r�=�!/	
���S��wM��,�~6I�ᡴ��ҁ,���-�O�o�C�ƶ�m����u%�d�C����@ݻC��.������ת-g��A}��l���˞��>���[%���i�Ԕ�<��M">�0I�3�d�H�;�Ҽ�i]�/(z��o+�)�������f}���/:���ԿZ��j��д.W񿑭�FJS�g�^�6���s�׳���u���<p9A/e�29�(����	�=s�+	�@�Q�K��t]K�H��Ϙi���������'+�;�
��������b�N�g �̱xH@h�d 	?�X.��u�/�ZY�Nv�[5��3��\.�R��)o�l�ە���r]�Ig_��K&�^=���O!	^�����bf�����1�ʡ$��5+����3����CA�V�����_���}_/����
N�
p�R�e�M\_��<-{&�{�i?�Ri��v�ŗ ����䉟��M��y��{�yS�+[�-<�{^_��s���>�]���]ۊV�j�O��􅱊 �Ɗ���QD����X�qC.&�r�9%�]�d���/��#>V-SY\KB�8��3(<n�a��pF��sR�:�V�j��޿;�������A��ܪ��jjU����\?R�m��S����J_92i0�J��J��7GV�Q-��}�zx9+���ZUo��k
1����>�{����e��1�6��G����ĥ��h��\6��h���`�G0\���N` %�<bD&���A�HuK��L���/v��ՠ��������3�݀R˟~�����i�m��taY���9�����Wv�^�)��\FhӿZ-����QC{\�ۻ��73�sg�k�/�5���2�8q'A�s2W���qL�PK��_�=��i�_��/��=�~$'H`�yP���p2��>8te��������^�.=?�\�m�ń���G�S>��
p[�\�&��)����7dg-����N��=\*�-7����Rx�6��1���X2`R餡��j��/��_�e~p�jSg������YA"
�n�檑?�r�]�P��=�'�#�N+編�MD��aeu;].��Bm�cj�>�dQE��ۭ����:�z��|U���h�rLGhh���%Vt��;Z��bM��1���+��--0r:�}���K$0B��珲Ij��m�C�igAعD��s�%u�D�!ÀE�ts�w�@��O�<��IyI��F�w��F�B��=��P%�k-��2��_��#��>8-�>��|*�����.��
��H�y�d����9�uu��G9=�_Jz���Hq
#�RMs{���t#�P6=�u�D���+�o�3 �{8���+�#��>��j�;x�d�O�|�H���	M��E��Ӂ��]`6B[�g}��?i?O�L#4O³+�a�ʑ���q?_y�zD�����r���,�� -�4�Fi��k�*Y)������H@ 3�Je3�������1�u���&Ht�d]pW�i����3��D������)!в^�~ɭ*�"���񽮗��e(-�b��}qj5���=t���2��L�z��-��Io��j��B���	�O&�4���,I_>-�󗺐�e��&ͅ�A%!��A�5���/����v��ј�ë��n��MR� ����-%»KO�����2�dDWNU�m���d�M�����R��q�5���w�f��3��P�*�M�f��<j��;��ʛ�h��z�lɠ*���F�|���3U�Oeԏ�;�#�����w�A-B�H�T�-���z�����F�Y�tG�*�K�3��P��/�w�)f[`�K�=f���H"�R�~B`�����&"�!�hXV�]9��Κpg��0�� �M4��g~~~�d:����
���D���x]8���RD�1sR���A������R������G0��Ԏ����U]W�T��[�_� �/v�3zS24:�&q9I$�]������5�@G4K�%����AT�ӯ&6Q�j�'*z�÷��N�zZ�>���^h�ŪRi�x�a�����}`(:�� �y�<[1���/Aq"�x?e����$<�]��'b^���>,�d���n��i
�R�������L�#��f���F��Q	�q!?��p.�`R���8IA_��2E�	�ZX	#��r� Ŀ}�uN����V����`M����GaI���|���/��okhե��3L�n���n���K��r�h?�@1�����T��v;**؄�öK״�ahi�\�D"����Sy�J�8jÐ�>[Ep<�9M�հ�`��Y)���N6!�19ap�!+ `�GR��y�����3ft|�/-�h����S��v���EQ�{��~zz���x������3PE�j�ujF��� ���v,ܖ��
{���Cz�a�-=(�b&Q� 9�|�Yͦk;��U�"g��&�+�kF��Oҗ6=ݪ����{�x��pC����:��2+g"��@��'�`$�0x��M�R����u%�E�d.��P��8 ���)ǥ
�ԡ��B-oɮ�~��y�?/��:�1�a�w#������я��i���D� P��e�S�tꏀguS�#!���B�LN�`7��=W��� �;�Y�xW����E���L�g�>�o	�K��"�&�ޚ�aR�����[�+[2����v䦓���k�"�!ѤJ.��g�C^Bw�t3��5��m�5pO�01j�+\�ɺ�Ҭ~Z�䞯�|�99�"���yn+/}��s�B$V��p��Y����.]�D���´��}��"���!бh�xo�w�P��ܱye8��i�\��������-zqu��f7j�~����z��WN�-���^#���&߹6SE}���:t�}	�ߛf�;J��x�9 ��W7R���
��Љ��	�aR�Uſ,�*"_k�����Yg6e<@)��W�Y*ô���W���_�2�n,�)��]LW_d�F<P��|o��L���C�9Ӄ�ڟ�x���.�A1�����Cx�|���4�Ӡ��-i5��^�Fɇ���J��o���p�4˔��c�xc����������5�N..3�"m܊��γ��:Ii�՛�D���^3�`j��-�$@��`�:�q��:�	�<��J`���h���K�5u�03��<4Ґ��*�y�㋗zsѴY�x��V0���C%8�������I���1�K��xy�+��r�f��5y]�ī�[S��Ds>��+��c�;U���` ��\(&N ��	��ך!��l�XjR��X#�I�iI��QN)"?��1���*Ř�v7��5��h�4�;I%�1��� �u�g�BA�ѵ)4l@�x�5jY�DSP�4'���[�<�--#FLy�T6��C��p�}~���o���)�8pc�8e$�?PP� c��L]�#��iJ����^�V�>L2�h9Ҝg1����g32ni�����ƫ�F�h��:���Aɔ�Q�ner)�\��S����z��a�c����E�Rʹ{Ⱥ����+�K�Ab}�
#WR�A{�l����	n]օ]aLv��1��X�v+�+T"s�P�"�}�|�5:�:N���Z���������ש�7�*�Fm�E�;���k�mfӭ_SL�	��
��',�W�T����p��{��=x·e�.jcث�ơ�K��WJ�ż��{?#�l�_~��6,Y��:$J�BpI�"J3S���X�����z���=�,{���\��Z�8��f�r�jH��mk�8�q��������Z=p~4zc	y���9�$Š9-��
�
7��}v��\�������T�'���B�K���6t(I}y� $u�1�V�c��I���:�t"�?)1_e����=C1�d(�n*c�2�;?��bkҀ���mteB9�O����$�ę�i�^ź(n���2�6r�Uɵf����<��}}�_\\������N_]�5�������1�3�ęrB,--�<z4}����W=:���bYڍ�F��F���p���<���T���k�O��{N���˳4%��C��z�������c4��3QT�Z�}��Ӻ%�>p����w�7�WXa,��U��Z�� � Y�P�${�X���!�q�s(|'�I���;�\iH����yJ���w�Ԯ9��{��xgݺ�K�ɑ� 9�0W<M��쭽�U\��gsC���dŹ�xzd޼������/�g�1w�LB\���]v��o�9�䍅�C[^*�J>n���]_}j}����+��P/�;��јGq��白��Ўa�M��Ÿ��{�!�mS:��J3ĉ���庿}�����Bg�FDk�h�Ud̓؂("���GR=�g�/��7�q�{y��n�/�%��M�|�o�Ó�=�ezj��z��C�ʀy]�����%��&?aQĮ��o�K�����=Q��f7�j*^��aD�j�J"����v��ؤ���H�N�TI�&S�ɡ�������͵oWY�YS[_[�C�"T��K��2� RQ�Ֆ�����C�agg��i24{q��y������EL�Y����Yh���M`Ą(7�WVW;<��l�^{����$�|�P���%���X�W�+ۜ��X�I��2���'�Zj�U�ߊL!��˹�È���0�y�BN}�?��u��7tY,�R8q�~����й�
�F@~yz�$�����A���W³/�*�f����g�cC�҇.��7�.	�g`����d��������Uɇ�3/ߋ�UԳ:cD�K�������L럗�����OI1F���O��b?���E>Ź��9,����u�� 	q�ʨA4� ��-���d��T�9���H�*'d����QMZ���5�ܧo��k����&4C�ؗ�l�%�i��r/����X_������x��Ga���y'g��$��t�J������N�u�L�BQ�?B�w#Z���N�WgjX�H #db�>���S�/o7N�c�l����FJ|�i�ޙ������!��i���&�̝;�C��_>\(�Α�F�����F0��x�[z���K�H�3�����Ӗg?��L�f�b����0!<�5Y���_�̐�x	&�8����k<b6`R@x \�@�L~9�l%t�9cꢻb�Cñ�~_ti$-{_>��O��;��� ��A ��G�ss	/��{�������	�	��lͳ�&�i��\f"�\�C�d�3��hoo���z��MLg}qA/��B��vf���3U�Y��}>�mL��;���o�|�ǝ��5�� ��k`�8r��H(�	AwQ'������;�B\k��t�s㚧7n͌�'?�	�ҿI��G�rɔ�.�R�������y��8�q��v'�Ր�G�4<�t�:�������L\��84mlV�H?�1�9C=7P4�&.�D]����i�C��_ok鵂�4O8N\0G4�L�,Q�7�̌�M�bT�&�m��a*���9H��*~G�HV�Y�zTI�Jt�[r-���D����4�t&tJc�R9K��T��dy2�>R�����-�GK��|�W��@돞f+���zl�hؾF!~��Haā[u���n�ý����*����,lX$��Ɗ&���j[g]]�?���A�s���g��vj/�6@ ������яn�����i��ip|��3���cȁ�Ϯy(+{��΃XP��2��T�l�+����j��i��^I� ��"g;E�n�!M�7�z+�L���(Gm�y"RZŵ�WΒx,FE�)"TĲ�K���;�-�;����̯q���17 ȅ[�������@�^3�vg+��.?֓��r��E��;���e/��:^��ґe���+�E����(2G����
�������=�@�a�c�����&ixަɧ�7� �](*�%�kU��h&�ӒQ�9��8�@x�
�ܿ��PE�#x1`�Z�7:\c�x_�:r6��g�9�H$�����9���C����@��<~��n�BίN��A�>=��z��Z�"Ec{��'?ns8����d��������و��=e�\�>3�K]
[!E�ׅԹ��,^B�4b�����g`��&����AU6z����U�f- �T�a�2"�{���H���N1���d�,�eU���K�صd���C��+�W��;�a����K�S]P0)-�r�J�f��r߁\ePA8���u�.�y�(B�<��<�_��=[�4`��0��J)���WZ��X��Y6P�~�1<>���@��X�zzb���j\�<�u�l�Z�JB���e�#��C���Ha�N`慇�:D���IVu��Y���:S%3�s���***��?�M�D�����Ŵ�(�!);�!
�Α|������P����F�7SQ7�0�+�e�L&���E�i�/�B��ԷՅ��U�x��=R�d�H��W|����Y��0�(����5��(پ�j9F���NH��L�8�q���I���N�b�v2o&٤��L^�R��qs�y�<u�g�
�`��5ŪX7ubIdea�<x<>�v�$����7�zlZ�j�Q���pn�s�3u����?^n�g�� � Z�G��}���B���7�o�V�2d���`"E�@�a��GNKKK��
��e��G����8�HſŒ�}����S�7�jFJ�&�h�
�^�6`����'p��R�(9�J�Tst\r�?��0�T�_:i�Z)���3����w7���}}.b|�²>,�a�:U�_��Ze�����QW9hh͵u��#I#3���)�<�9Y�bH8�{o�I«<ټ.p��^�3_�؄8^4V�<��a�T�Db���/+��v$-�N!THY|��ٴ}�[����[�?%0�0�'I�
{$9�\�L7��fG9Yv	q�~}`��RAi�4�̵r�������S���圹�F�!�y�iR�E�f�]w��
jqs��@����:M��F�L��t�����\(�����׍��m��P:���n�Ϗ���:�7�/CN���(�a�Hs��b�z���h��׆�1�7PM�W6��:�c�#�h���̕�wz��	KB�}�r��0�W0�D��O���{ �Rkĸ�),��i����,G� 4�DvJ(-�t��3ڶնAY��%,�?�נ4�H.�ٵPh�:K\Q6��U`HLܿ ��v��
���P�?>��>� � 6�Q�����A�5M��L��Ӷm۶m۶m۶m۶m���=��_�3�V^��"J�&6�J�H�'�G���D	o,+��5f���`�G_e#���o?�S%�Ӣs���{�ƙ{�g���RI[V�@���J���V�l�})殳ϕ��{�hPP�m`v>>tI�1Q^��O�A�}�������i��rZ���4dz�/�wh�O.0mwyp�?�<��aƑ*�6K��/6zB3e�P�z�����B�b��B�4�I^#ڲ�����w�=�q�-AUY��>�q�� mB�5O�/T4T��MMG�Q=4��h�}@J̖b!�&΄2=� ���$�}��#�1!'ݖ�U9AJ�BU��/�_�H-l�/����_��м±E� ������}����Œ�4�eײc�u�`KM�O}��oX8Z)�8�b�=��i��6�Œ4��Êg�&:\�&ypd-e�E�뼑�>�F����xGp{Co���m��g
�'�=�Z�"Ig�#�C��̻w9%����5��6:�Lq�����y-�)���ic1�e�����L��Ps(��Y��ӈ�Pɨ�'�{45Q�+��2��?E
���ok���(qQ�l������cG��o�\�p3�]I����<>�|�Ƚ��؁��,f�O�l���������o� �����������}�(�2H�&���AЯN'�鏱]�{D�Cr�W�X�zE��_6�l���SM�99o��ec5mN��i���΅�����sк�7$s.A~$x�cd:u�V�9�"༯e�����
��T\�nZ�f{d�ios����y��X2Mm0؀��B�p�4�?�,��|��;�a���w ?bIJkYU���댂�2��ci�RYy8�5833�+�U��-�������V��%fK����涪��4<��c��@ժ��;1c)�}�g�$����j���}��S��&������6��g�}�e����W���k�S��f��-]u����hu���c���j��r�󥇪f��2��B��F_GbT�tN��+�4Q����gO�צ~%X�b^�8�Թ����g���Z�!��㎹�6��s&C�t�[N���ɪ=���C�K���ײ��ЧZz���s��n��7�^�V���D-U_$G��E2o���`��<"�EK̱�quTK���SR���YQ��t�f�#d��p�<&O�r�{?�g#�m`Ÿ_1}��ߎ��?,��Z�5"<���H�1�{��"���6X�xs�^[�lV<\�Lu��C\�~B�ő���h��X�k����O�	�{�H����$F�!m�R	����C��/�`��b�O<3�X/�UNlP�tv]U̘q���{6\%kx�g�R�j�;\R~�z
S�Њ�)}�!�A��W�WT�Vl��$��-UGW^��q�I����ի�5iqKv��H���jKKL�a#z~�B6W��\�d�{F3N��S� �5B�r�0�J指�$�b���з����!�O��S�Ȏ�yɀ���y��M��>���ܝ�8U�n�I��2��Ѐ�X����Ε�����>�w�h�t��Eeƈ�h^����=����u�����Ƙ"l�+Yq斍0��Nl������7a���}��iiv���� `eb�zU�E��e�;@h��*4 ���W��JX��:���m��(I�o�֥�6��ؘ�,Ӑ�E�"� �E��/c|���3
���ٗ��"\7oW��n)	�2��ys�F̟S@xa�����C;t��v��D�9)�j��2Q4�xL�nh��U.����Q%���\�'��8.-kR�/oO��T��1o�����q��\��
�n��@�l,�L���YHm�
��u^���k yw�9�]��j�J0ŴG���'�g���RK�V�/�|�	t��o
H���k�j0	g��N��g6#O|��4K�4�}��cG����0������w_����:�������1� ����������C&���CfV�{�����fH[���J�������J��qK���/�Ga��W��|[T�A��`�����̙2^����k��H�S�,,RUы��WI��5OMe�����2?�ҕ�q�@�C|��K&:��#w����6���)f�����3?k�/EHa����\aI�q?�{�3��tP�u�EYe�mjPoNa]���z C{é��y)�Rws�y�.׀�w$�RAG���?�fڈh��A�|�ܕ�hmC#��l��=�����u.��e�'�6�
J�d0����jP�n���;�`k�J���ńV|�/����!"֨�p��ddd|f�����������ti�h�,X6�fX�Y2���Mʵ��û�Q��iՙ��{�i�~ڶ��D,']`a^u}�Ź+ə�y
�����E�Be��#H.�l4F8��VY�	i����,xcr�t�Ѩ0!��"��`��6]BE�}/��IQ�IKHՕ:zNNI�B��R���X���{�����R�)�	�c�Ne�b�q�P���/�(aB3yq�aYq���#�b��xߥ�'�$щ�[NX��(Dt��XB�3��9+�4�wU��j�P[\o�H�H��{��0��zq�;P����5V���49W���͐�
�Ξ^�1��RԼH��:�B�;�6��zuc7�"NX?�<1����TTl�X@S`P)�F`Sr�P�`�s�/�u==1p��tQA�N��qJ8 ��ǳ'��嫞�����\q$,a�r�8p���!>hA,
-:��3n�M��A��{���By�8�p�Y�s���4}s3NCC�Dϊ-���g���66GG��*�ћb�\�r�y`��gtb`���=�AQ�f�5�H��I}4@�g�}g%˹��i?~ůg����Z.U&���Ĕ�����Q�R�)����6�+�8NB��Kv�g��"sak�UL]�7�����q8�i��I����7T� �"��P�c��U��Q���i(�\�Pu�A��sI✤Ԝx����/�}�� kN*z%������5J�����J����х��[[fP�B�⾈�>�j#$��� -Z�C�reY�  ��"iZf�w��F���1	U��bdff������O��4礕��������4$�k\�̝,�P��:����C�vxr������4[���&,�'d��>R���F��樂,F���׬�l�X~p}��xO��x��mSǴ`/X�����rf�[x�0�23��FL+�����I�X��;�6���-r�����-7���67�����Z���O۲��7�	��+�<�o��������?`~�ᎍ!g��q^�I��t��B�#�gA��ƣ�#PJ|�~�)����v��,;4�eON�|�Jܓ��x
�Pj�^�wH.>�}��#s�\x�.�x4��x�J9�"����b̜�O�
R.:�fwL�̽�!��@M��$ʵ26�'�����P���w�x��V�+}u1�۞;9���``���GIdj�J�����$�,	�XD������!7\e�w� dGcB�����h(������of�\G��;����R�LZ�Å���s�^����b�
2E���?�0e�`�&O���.�U�Uʖ�/���#1


ƌ�37��Lg=7-:;^6�8G��S)���9���ݟ�u�^hs���u|G¦d�D�ܨ��@YR�݆S�����&�� Fd�Z]�U���;"'��^!29��'�)��+F>K	#-�����@[ӥRBǕ+ʷR��Rr��!<�1Y�uM9���h'K��sQ�b�c�	a$�x!1�ϰ�ՄN|y�EJ�d� <p��z9{-P��O�� ��l1C�5#�K��L�ge
7CC�O�n�z�̛�l�uX�.�oܱ�S9e._s�0I.�/<���c l xr��2U_G�4��Ya�<cT���l��ti��v�8@9����nb�{m|�Ju't��CZ(R(an�)s�ӳyO����9�I/$�F� =�Ý�aG_�v�K�.b��hkGex>`��b/�����T����V�*A���h��r�m��S¹�q5�B�U��A�1�{#�e\�W�Bk�J,���MQ��S����llR\�]��@F;��"�Kc�p�j���s�@��R�ټ��g˜���MN��+-R#���ؓ
k5!����a��p�SxҸ�n�	���R�r=�ϼ=]ϼ5��`���}�pym{f���H�)$�a}vc�幐IyYq�H��[-Ջ�1��@�@��^]�UK��/d�F���(��ȏ-ʵQp�0��m���m��zݱC(Š��p樭n�#5?����D�	5�f1���,?Z�/zp�~���&ϴ�� �C�����0��a�7�&�p�[�E�|�]�q��Y��{�����X*!�E�/�QH��y��m��ѽ���D��f���e��c�Fey���@O�D�D�e
�r`��y��E�����	:+�"��MY�͟����i���,�&�0���=S�ϟd0(nB�d��Һ�+��m#3uQ���I��qr���3��l�B{��<������όg@�*];�Qtl�>���m�k�o���Y���%���O1�bj�%TQ̗�c���7@��#��%q�����64�U��G����[�yװ���փP�_��J�(���Z�?�f����V��d�~�#3�;�2d�4�:�m���TKɮ6O�;�9�o�^Y�	��
��E��&O��36*��/��|��|��B��~����{��������������;7W�%==`��^h�Ufϊ�r��tY�)��e�<S{�n֜�*Q�Z�ı K��D쑷�SJ�}ϔp��ʋ J�����w�g5i�-����<-����޷(<�\��ʭv z�vvaMOL�I�I�F�
s=3�o
�~��;���> ��uc��CbmB}W4���T��-�������247�	Y��V9*j����D���,�@�U��7���B�=��Xz9�{��+u��$��BE�E��޲ʩ��X�dG�3v੕�_�:�7�L���<�n1��90��3ʫK�S��4���s;z���]���C�j{W��VKG��V��ȸRdr�5�$�<��sx/�\�%h;��8U_x**m�._i+�G�Ӵl��|�$ÔAp!��a:N��(�z5K�;��F��L<�hdQ�D�f�`�j����֖�e�Hv(�T��H�,�Q(�''�6�%07����j�����J�Ya�
�:S���i��:�@39TR�H	�l��SY�Lj�>r|�X�MA����m��m��U�s���+K�e��9�L���+ؤW6�60:A�a�q�KP�.��)%�L"��-� r���*�rTT��������;��q�hD�Q�����8jb�����\��<�0�}�}j���d�ȣ
J��!�`��?�dxC#=���Bvn/n�pR���k�8����v4��"-��^�^M���;���j`P�����9�Ի�s�v��XB�F��6���s-"S �c�ɩ)����Fh�c/2	���}͗���$������j��!,G�q��g�������Xה��Г�
�B�[&liQk��~�D�փ<B'��p�IhD-��R�A����]f%Q��ۄ�y6�8Av&Y��p��%F�59��Ab0A1QIY�[������������8��c�C�����ԓ����y<�P7��@X��ϘKU�MVW}x��m)C��	l�н����{�m_&M
�ċgίsJN���_F<�=�����ۇY�����GM������\"eǻ��l*�of�b'}�_E���ߋ{/O�W����"��ƍ��n
`8|;�O��}
����Q��%^�3tf��R��/�@���>����éޟN�m�WA	$�WVW��%�, �!�����ܓ��y4.?~|�u�If�����Q�={�Ӵ�(�=8J�4�e�+��)�,�b�^=�Z�h9Ǘ�����bo͎ "t�U��9/p�h�)�)L�}ksk�ԋRnjX:�ڰ�{8���HW�`�>k��z�Z0���9�:�:���4�(L4t�M+P�����	~yM�R`��V����~fZ@˺�#BF~��
�5t���$�K�+'w=>3��'���t/I&+$�5h� GlC�y	�F+wD�]�6`��)�rN�����=���6��Y��-�ڄ|�Ź:��UpÉ�@��Co2�bO/^���O
dB�$E���qEGl���`x�0��/�R2�/�&ІB|q'�w�E��!���dH��o��dLK��$�2����R�����\i�Ѡ��p5��P
��mE3ER��d���iU��5���"2V�뻛��ԍ�������Q���XTut|�<��\���v��*Ư�3<+���}�n���$Ӱ�-*�l̾j>�I�4`Y��^��C(�!�%�is���hF=ǋ��uu
���͌U|~4P�bsæ�;]��X��a�-JQ>X�3���N�D׊�x���B�Q�A�:�rJ�C�<i@U_̛7�2�/����׍5p}܉�	�'�����M�ڝ	!�D
 \P��C�1��9��6Z�df$�?z|!4 � V��5R�;g\�F��`^>�]������S<o�m�}S��Xϛ7��}�\\\��̕!l�kj	�+*J�̡ȫ�_s��f��Cy��ae_[P5�������)A�s�88{����!����
���;/	T�Ȧ�l�8;�������=~��{����;N#QN!I�(�+?�Y��>��FR�Vc��=�
)���.�����c/��O&��{4��x����}���&�u�K�h�Lp]@���E�k)��mb�LF�g,84=��e�Al/���������i@f�X�n��U���wO���$�Ӳ^�!8t����c�9��{tA,ǅC��W�Oo��W-$:3�aw�⊟��$ߕ t=��D�}�����L�"�p�1���dW9��U�#PWR~dҾα�%#X�T����ڶQ�� g'�5-6�(���}��Z`-�.�_q$;2�	�튝�Bѵ0��<J�q�T��4�e��������P�&3O9Q����-K��ud�L���%X� ���륹l��s��@1	�B��l|���Lwm�L�u�z�����I��`b����̽#��'$�n?l;��D?t\���:�q�V�:�C��Z�z}*�q�t�W'9D��T�WϬQ��<r$�>$j��z�{:9�K�p��c�J����=��^� ����������q^�C^�#�l���w+�\����ؐ�����]la��x�1�i]ȅ���x�����U��Y�ʡ�@r·�pD6����]�ۆ�vK�C0����qG�q�h����=���ǰ��-�1�Ё���j#�b �S)���mHR%ZT(0�j/f"�7�H<)�}�n����Bb"��eק��1�a���R�:�@zC�i��������.~	���#���Oϭз\2�z*�=0���0Pv�y�ns�s4ZT��:�����ut�5�g۔�����]5�1�v�R��lC�����l�NH�� u,��:�+;��K�%��\͡mۘ��pT�����8�aU�`�bb/��xd�8�K���	�:�d�������R�'/���&l,n����/~��VU�pA`#x�X�������p��9"�����j�x�����6�O�B�P��A�]��Vʍ�V�UR����$*�!��Cͻ�шL6������.Y�����I�3B1zH����|�b��&u�d �1����������(!)�0AA��r�2�5���N��6�,mG���/��Stf5���֓� �.v?t��m

ү���D)�+��C:fOl��;��w� Q�l�E���A���`@B���i�bf�yӯ+٢��Ԧ�jX���2`ʤ��s�+9��Ì�>4<<S�s���\LA=M��s�yV���u�����TLp�2aDG�r�2n����ee�Uh�)�89���3J"2	CZ5����6�l�X�$�=�
^����9��D��E�ܐ r�M>jU�!Tb|���盜Z� _U�ʄ�	�w�$�������2�]�h�Zή�H����RTg�1<2�v����i�!�p� ;�y�0���42;�$�`���u�j��?�֘0��mڌ*ԝ;�Hͼ����Ǯb��o
#t�V%��1�@�ޗ	v�^�^<�;zG�84~=�C<���	i'��<�"G�j`��O����y#���⊮��-��a�`	��W>��W(!/=�f;=�b����C`��BF$dg���y�)�h'\��:��|��΁�;8���1��#�p�ߧ\���>4$.�)�-�l���$��JX"�8���*��| ���r���1��44�+�ޱ�W���8��y�ZFV;���i���,��*��a���8	&�%�T� j��V7mO�W0T��@,�]ı��J�'�X!i�+~2��;��w�3&�3�ᨁ#���X}���r��fC��{���s����C��@�ބ�Y���s>������YŰ����>���1���2ӊ�{��s��s��X��}����c_4ܷ'������#��T$5P�Pj��ޜ�zVՠx��٪����Ǻ�`�ѧN^�^KU��������&L3�j5Ԍ���{��e�p���yt�� �O�Z'�6�St�)YS�oR�E~�>�Q�[^�da�� $�������TV4��ח6��_���
��������4��."PƄ�辫iQa]��#7nUd�ag����l�D8�6p_�c�ch�d�ö�����[������:&�����@�{F�[��Gy���[��yƺ�Hoc-����DNrP� ỏ�|�~�Z���
��U��;�}:�O�<?�j]� Ą���ȁ�uxc��"µY����A���H&�l�q�oy�.;y�0]��P7��9�q:%0,�*�0 _�T� �y�>��_smm|���h� !�sPˉ�݈��Q�0Ҿ� ��=�A*�V��Α�E�HO��_�S�Gy�<�*���Zm�,n߰��-o5۟�����=��^�yk-���.O��*�������� �|��)��}4�=�Y{�����,έ3�}@���,��l�.������b	��|���r.S����c�}&�N@4֐c�ދG�������eI��ƤG��	HN��|A� ��$��U:-E���B�a�4-�sO.I�A�,�>q>Tޜ.Ac�<�M<�k�q�T+W�ox�4�R˿q��$��)X��;���HCS��z�ؠu,+��#R��ݥ?nU	%Op�Ev��\�C�!S�Z�BJ=�De,��NX�p,�H�Q�d2�<3�0>s��:Ň�<Ë�_��R�u�hl[�=��,��?����l��$9��X�����Z�\�2d���V��&c��b���KQn�^Ng�f!��n9�d�D���o��GXC���[��C�������*�׽��p�m��=�S�SC�Z(�D����$�TH����f���Oأ�Ip��Eׂ;���7/��X�`�^����������Í�!��ck0��p�I�Shi{M�]�8+`����b�i�8Q��}*�Z����<!4�˕L�;�����0��XǼ7�;�*+߄���i«�Cb��yAC�L3T'R�UFȃ �
/�$��x~`�A_����RnZņ�e���f�uj�"��H��0P�JF,�~%�gr��cpJc�-F��r_�1mZT��ڨ�������X��hI��P�%q�����	��wJӞd, !��D(z7�M���o�/�hV��!3]c�t�?�Ŕ��\�ԡ!����+��w�A�� |����p@��xc�f'���g�'���{�vf#'n�	�&+�]l���bb��k�rj��[�{`��ӑ#�vmV�)��d���=%��
v$�F�V��;ƀ�+�����0�7sFJ��� <�/_��ˁ�Iz�i��v�	Ek*�}dA�q�i������i	��B Ƽ3���X͏�C�a�h��^Kh!���H,��`�X��B�s�Bj�X*?����Aq�`�]^��X
7�g�������{�W�>ˁv�D����*�!U��K�K��2��������Ҹ(�٩W���8�&�x����C�,�{'e��V)�nt�b�%�/�('���GrčR��ѣS�� "�#����[�|������xB:���j��ʠ	>��s��ެ��)0�R����fka@��c�nhx�"�n�!([�?p��Y�~�q;(#DXЍOǗ�E%� ��۪�HV˻��^��5 �k�[r)Y�M�jd��� �qA����.��N�EB��5'�l870X�住�FԊ5���P�#H�x�R6;?������1���/�̃�T�^㲡�x���ң�5��7U����>�a��_/�C���ˈP<�!��ӂQ)icy����迴���%>Rk�T-��!�0�	�Ϝ�r(��狿F�5��!0H"��`�΁�mKv\q�:i�BA6u?P"�>\Tȳ�%d�Ud�/W�l�06�4d�m9V0t�k��U"an;��t��l��Zk�[jEn�t��S����̋f`��$ǈ�~<>U��%�>1�@̏Yh�5M6����2��.��l1�mE�'��9�Y�$M5>:ʿ���͢X��4�8�����@,ɼ����uSa7AK'�!��,j6�0��1�!B�<8���e@8�Ϯ�8y]HH�C�-yJ������`Pp-v���P��\�7ֲ�?qs��v6V���@Z�}�y��r�=���\s ��x�TE=g�V�	r��Ɍ�}���B5��0h�W_�	��NSfD���W��0��Q
�r��<�25"(%�`B0���uv�&��%���d���!Jv�;�g��s��S�t/�vN���t_�.� �,L�7Ǹ��[c���UWZ�5^�{	c�̕�����
��-ǉ��+�	�j���&�}2�BL�q�	`���b�7��+��,ռw�Q�11H0XFn�3Z�؉eG�$������{�d�ǽz���1X�m�1�*���0_,?oӷ�mV�}�k%�S�����?<�;u�Ib� �\szUS;���m�V\c�X����:�UW9ec���6-����S��n�>1I���:�� ��*���uۚò��]���N��.�WGޖS���}0W�/��&���n�S��ࢆ�NR��s�E�E�,E0�e8�2��~��x�x|�����4o�b��,����ڷG%�53������P�jL|V�|�|�Z��`q��}�*��,���k�K�cFG�cVחv�?��e���\H.��Hi��0�h��(�>8�>ԒPa~�����k2�I��ށۋ�]�7��-��aw��ꄊy	�k� o�����#�1�y�����B^��v�a��=�5���k��SsoO�[�BX�u~��[Yo�4���=iwTH�V�]���۶�;O��L�lXp���U�&��a"<�z�h��ގh��32Pd;�sD��FּwZ7Gd�a���{T�s�5��>���	q0~�*$��
�!H��K#�2��n3aQ�� �)�W=!wƾ+��a�P�m�?O����=%[���qձS�6��{�qSjE��EGc���E'N-�桷M�~dT�w�\��<�X�����q,�8���ZRϟ&m]�V��0T��j���Tx	z���u�)c�%�LM������CTB�&4��i��et%�y�8�~��W$ω!�!m[����G~0�w�2e8?)m�zJ�)������7-l�#ɣ�w��`>�G�Zc���#��5��b��>�+���s���s+��R��\��e\A�t��g����#���n���/o��p��j�1�=�#�3^�\�2{�""��j2���ϒ',K���!�M"%pQ�~}�8X��'[���K�����z)D��^j�F�+�R;.��x=����K���r�J�	�����h�|:W�f�-�~���ʚ�#�a���,�A,w�Z��%<�!�L��k��F�%+��TT�R�d��w��
����
w��L����%�E��B6�&/n j���Ұ.)騬�S����Q�����8Q��⷟����m�󩯞:5lWl��q�kBW%�V-:��I�6��q���������S�w�z�����y���+�iP���4�(�Z�p �0*�t�)��"Ϡt�f���L�~��]a ',���+�+_mh�x��NEψO�-	epеJ?ʧ�W쇲�;4w���
&Pr	Yֵ���!(�#�ӵ�����S��Ole�k�OG�k� ��T;�"��v��2$���d���Z�.���na"u2�<��B�
5�4��s�P��I*���д�SX-��3 �nNg����Ֆ����������p��� �*f�b�a�a�!����*�V̖NΗ[%��*���c�R��R��}�xa��x<	<�m��L��u�=�!�J�_ 7��̆�m���Gm3hg_�9����\/̘�5l�(�)�c�����۽�"8w$)?�����D�}n�
��]*_3w�(g�dܝ�x?��<&&v!���4,oG�ߞnA������[�5��
�v�{󰡫�'/�s,dGt8�G����M�F�+�Q���2�-5#l9��B���[�?"��NXw!<G���bP��3#(��_d(��3�/�u59@��Up#���(,R���b�oEf㺴����J��ŲJ�����tC��є��c��,hexB��S��kb�p:��
�9)�A�;{~jه������^�G�p����c�}}H�Yl�$���� �)�+�gL���.���H�P~Ϸ9�
��%�FIT��8���F���~�w�a��KIL����t����D!��R�����&W�H;�ڄԤ�L''qւۭ�R+DX����=j�q��M���2S�G�I�'�͛��l�"t�*�'&�"2o+����n9��0�����Ӻ��ҫ\#�S^�G�ì�£-E6,h\�7wE�j�M7Gz�Q �	��w�-�+��?��_�yO��p�Ƕ�׶@5T�g���ؤУ*^zd���\�Ї��{G��b�'�5q]7�&��0h^Ќ�ʤ�F�J��d�(rD��G6T��+�27"��c��
�RYc*<�|���w�jFl�+S6����,�bP��oG.{�x��{���g^���G>\6/����n��A�rÞ4�9��|R�r�}z�b��1i�{&V����^uh�x%hn�>�k�űq:�
��P.vvߤ��JwHH�,��e�����'H#��<v�25���[�7� ��k#Z�Ւ	��kV2(��_�i�pt�0
�ѢC�E����tSǔ�2noS>������u�?<1wA��4k�������V̄�X��CUʶ�5ft�+�����>ng�5ha�
]��y��E˨^����\{��Y*��{p΀-Ϋ�}a ������51=)'?V�0��t��L	C�$���R�.�\�ư���}Jd�|/[��w���{A�O��Y]+�S����Mv 5�[xԋ��W�;!!!/�L%k��8m��|�궭@�6�+��:H�4���Er��l*�v�fQ8U��H�l(�� <ң�<���E�aC��U�|��Q���!��t���^6e��&�(�S�"X�������;��Z(�	�wu����tQB��}��|%�F<����	J�olU�B��t�Rbf�f1{���FK�]�����A�ׇ.���� ɍ�ҶNpg�{�蒭*�$S]}^�N��,�n����fԮipHv�	�Ⱦ,l�{��i�M��ZF���Rt()��A(�*Jv�"�,��@����L$A�t5�h����+�Mb�����O��J�Kʕ�;v�H��^��$I��]-;��v�Z�V�=��i�ؙ6�����F\�E
�����y�{�"��`�0�` �3��5��so�CΈ|]�D-�2����AU&�����C��c6Ap�+�Y�5@qDNQٽN�Sw�u�����d6��4G�9Qb�Je�CRz��Th��7=������oj�Vp �Ec=F0tqI�-̡�ͣ
*	`������w-��5���c��S������6,�]��iJzh�9�R6��3)4���\ǌ�CtP��<5�l�C ��5�C���񺃤��b�{ݙ���[�d�rD_�,�Q�W��O	��+쑲l��0��и:{�fn#Q�Z���3(�P��]�����I��<��$Q���Aa���Y�%l�؃y��!E� �=���sۤ�>����2�]��4�/P�]؟)Vߖ�+���F��!��6��{2?n�t���͗����ܱ��H��;�52��p�^�mv������'�,\��I%ώ�bQ�t��/n�����c�PE�R~I3SP,궔�12Kis}�{a����k{q�Y
�Avb&p����M��_]PZ�׼�פ�9�պ�%'UT.��t,�^�"$����|��b����`���n�Ќ��3U�J]���f)���+pT�M���DR"�E��^׏*�e\����}�>�q%0�W��g�QA�D��g�RXtB!gÓ{�\����g��]�~q��\c&5l���Br4vA^����\�ċ�X	ĕ�6�zJb��Ё-̑8���U�Tr1�>���?Ъ򫎷w�3��@�H��0�曀:�ڸno�n�e6�8/,������9��:b�H^� �a�W�4J(��YA,�������R�MZ6�&���8�9����.�te�=8����Ŭ�[p�R�'���j1�����
%���!�y�!ـˤI���t
<
��ޅ��Ӧ�-�:O�ؐ�ڸ�q�W6GKac�ۭ}o:��|��%<v _�q��R)=��+��<I��`�z�эRf��ܡ�ͥ�p����bk��ά*���9G<�A����&BEI��^'����w�e�{�����-�͡��.f��Ǔ�i������H�V�	l���_�H�K�7iJs+ G�E^�
\�8�;���S%�8e�l]�	��H��q�J��qp��ҝ$����4߬��c���(���]�x]X���r��%_� j��*���]��r������L�c6L���êW��O!v�}z��+^�R�����n�,Y�$�P����-9/�6W��S5Y�ᕣ �*؂�H�o|[6��^��ԭh�g���Q��@��a�\�?>]FV;��3���t����9��QE��jg�/HR6Fg�d46u�"Q�q� C�����U��;q}���OD�d�x@��PG,��H��c�?OM<����Zm)�@S����W�jt��ҢH��rJ�ЌXu1r�	�Z�r����U!�d�c��V�}� ��W����3�k��.�僭$�|ۅ���������o�+�m:���G������RhE���Յ�Y
���,�DZN�EɃI��5���n�(I���zҫ��j�	�8~��}��]�mn��H�^�NF�݆��p�XVr������)D�����.�^�be�ϖ�y��S=ʧȬ����p��#A�LI:FM<���y�J-��p2c�(w��1-��q����i��sg�&E]
��b�
�ſ"�'����e$c��&�����]��zp�Õ����?%�[l�慇���)E�c �E�3��=� 󜍉ڶ�-��_�]q��7KǈԃR�����V�y�����]�H$��i�jBe�yz���Z~L��M�v�`I�{"�T9s�h�yW�[s�,	�\�k�Y��|`���!�έ�	�-Z�@@�����]*���y}TI\�fW8YH}(IDcB"��Ni:�"�֟?������#M�;\�"vKZ}�ń�H�,,,'�U�n0jv�lF�nM/1�ԏ�È:iW�X��l1�5e�չR��.�"*2+�] T�r�5��?M�����g���2Gw��³Ţ���z9�U}��m��LG�%�'�[f�\�9��t����l~��z$M�=0<�?��́ڢ��e.`9�J��g� R%�MD�qӘ�"�6���g�����p��iR Gs��5�'��_��xs�!n�t:J��`����]-��y`��o�ٰ8�ԙ%�¨khU{/T,�_�U�״U���I�nXBQ:Y���a�X��S�A@��\t��.���kYz�zy��y����·�a�7�\�3g��W5bh����J�U�v�F#+��"�&T�n�.�uk`z��11�L�^�>�W�2тwI�	�}��0�7�b����e��}�[o����g�!wo�Y������/m�.RTA�5�Ӽ��UoK�4u��,��s����v��$�s���98��U]��L�~R������cY������R�:��B�Ugv���T�� ���❟�9���(�c��.g&)8Xj�f��UWd�s���ʇ�U��{#��	|�\��=�%�^:��|AM�B�
��y��f�9��	�}�#$��@���/�̥vV_ũ�?�q
���ܦIH��7�w�^l��H
6ڱ���0��Ղ����F��V���Z�!�&��"�gE�ϊ���b�+�|��I��־�h3���鶑͖�^�ŰJ�N��遘n��o}��-d�iձ�+^�g�����E���jqQa���8b���WAΘ����/]LR�21�gt1
��*�k_�����4�a��Sꫩ5�vCt#g�k��Z��\�J�It%J�.��	D�U�ʦW���13�5H�$��X�p"a3f?�w$bk��^�Íd�~/��L��~8��)����
Mo+�|�1�"�k�Nu^�o=רA
ғ�i[e��������8l��ݷ���b��	_�|��9n]�$�rv�Ϊ���T������o �ƞ�Ɏ��֪��'�ãm���yl\Ch�,ϐ֍��y�xZ�ٜݢM+P79� ��]�q8� 8 �;摰�5;b�]\��g�8֍`�*�iI��CW���{���'��{�U�k:��=[U��,�/��b�|2;�x��*�%�(���XA$��J{s��r����M����b���/rⷮMi������MO/<gD��[�ZuU3`��S�>,��>�욢._�T�8�ǝo�nƬ�]�����]٭�*ͥ���E1=N&/�Wjn8 ;�8��a�Ou+��\A[�y�����3 �Z�t|I_�:�xm�`{�8aƀU_�6d���+�x����P^���;�ev����7k��Ko�q������.�zu�N���S*�"�S��ϭz(�1P[�}z�r���'��G1`���ˋ�V�ͨ���4�>�(�d��R;,!X<�6N�Ֆ(�m��g�����k2�JLӯ�B 9��"������?2�d�=Y��2�=0�h�{��.i*�i�4������ �/�� ���z�L b�l�z�>E�31-�A���[���"V�\����Ҿ���%h��%Deϒ��v��P��&�w���j�[�ٵ.O0P��?a)Ņl�W�N,�W�4�
�ţ%V�����L�_��>�&��@r!Ȫ1^G��uʘg���5�ռ %k!�`}/�e=��-hWH�S�F�x6��UUv]3sU�;���!t����yNj�U �s���(��(aI2���E&�}a��4�7:Mu�@4R7Eq`���0Z�`�ݥ^�GA�=�N:?�f���\H��I?�y(��{� ��&�+1��q>������F\�F��Ž�2ñ��<���t&��
��'���#�Z,r�-i�`���N����M؉�C6<�
j��NLR���x�J'��q�ԩM���V��5��Ĭh7yl�gk��Y��d����gu� �T?R1�Y���{�V(�MFb�y�(�NQ`������>��γ*���66��M�F՝�F"�I\��M1���p�W�'m�9�t��$�(�x=2M���s"Hu"�\[����.�|�7���"�Y���~F)�td%W :l��T[c#Lmȝ6c�T��m���]��EMg���I��������n��^g:c�%e��"�zt���r�/��7�?�ع�O��2�!�z���S���I%b8���旪� =2a^vD�4�ڐ_�:��x'��a9����]k�@��������>7j��_�}���<~�Qd�KO0�V\��M)��m�h����i�������~���flVӡ��t��������B�J�.�h~�r19�c�؆/��P�k�>��XV�c�&񍛰���oa�BD���0]�L�yo�eKz�K���x|o�#��k�=�
sq�Nd%#H��k��^���{�ѯ'n���4فS���kBG�N�`�ťm�\>2�o-:��4KgA,%�YY4o�m�����_�����DS)��\%�TcUf
u�<�pn��,��E͓�'�%|ZQR[�x�(;��F�`vU}�.�k���YG�R�~��D�9�L_3���@�"��e���tՑ���Nza�}r���)��1���h���R|(�M��^��U��b@d���^&�o�(�6=�=E5��yt�Z�*���9�	�� ���-X�ڃS��K�P�?�J�vol2�tǙ�a�nG�S`����)˰K"Pr)p��|b"t>R��5�V��Ƕ�7K�����*���~_ց�u�|r��;+��Ѫ�n�h�����:��b��f���m�A���E��n,Mb/w,K
�?��*Y�_=ok�J)U��[UX3e��_~��Oe+�t�.+�H�ʹ�>�+�V�7�����YF(3zsS��2�dY���i�f������;�Y}ZNp��u$�����0�IZ<F��)���30i$>U��h�&O�U�����%���f�CD*�0���$ov$�Mu��%�/|��K�$�8Q�
 p�o}�i�>�X�����Uqo�W~[-������K�k��D�������B<��@�:�G����^o`�w��C=s��>o���Z�yf�*�Q��{��Y3�U�` 9=SwnVCq��F�R��!mǖLNxt�~�̽:1K�%Î���\tj6{�G�̬M�|��6�L����x|�N2UP�M��nJ���lz��/G �kC�-� H��5^*@��ó^���X;9��KMu�����ͩv��s�g��S���Wv�C>�_,� ���w��
�IUX悢����$�-v��ĸE�D���Ȼ3qE	�R.h��d�rS PC���g7<�R�~�Y���jRA���+�m��_;䶪�<L41M���hM�$����e$�l�^�������Xj��y �����h-��Ȅ'n򫟂�*$3�ϵ�^O������i�Xgw� ��4���)�bNq������o��ՠ�D9P&��۝��;��j+���>ø�!k�[C�fY�	��������h�����N��\��g�C�Kl'�����r����q/�Uu/N�;_���%b����wcJz����
k�^���KZ RE�fH�)��> �&�Q�?�ιky�N���������+�&�^3���y��*�rs<��u�s�i���:5���x���KY���+Q5����U��[P���"�T��y���t9�_�h�.Պ�sS�P�p��x	��O^9ſ����o�1Qw%���?�Nu�q���y�t.���9��Bf6��uE\G�fG2���|�����{=����HD=��ru��LM<�q4���:�}S���w��/]�T_�@�Z.<u�GA|v���tB]��8�=1���Szt�0�(
���C�5�黂�f��~�Éڴ#�w��3g����{�̟xyJ���5�o�<]�i�~r|H�	q���B���ΐw1C�B{Th�	f&��g��i%�ҧ[��I_J�k���ƍ�
!'4Ӹ|�L>��ıw��m>f�ݗYfʽr���W�go��Қa�Mb`�VS�܀7�����w�����#��R���L��O��<Hy�<t\/5~�,~]�М���0�*W*)�G{$N:T�g�^��M�GGE:k7�~�������D�Pu��=�ۃ�{��V�p6���m�%I-;͍���Z�y�]r/Qކ��Q�����,*ןf�r��W�02K[+L����T
�v|q5|;m�'{E�+)f]y$��Ђ��(�6wΏ���ʴ8N
��5�1KOy'�jʖ�S�dGk�5judt��ӆ��9�]E��<����]���Gx���'�n/��v��4�1��J�������htLj��	G|q���:�ɨ����oB%W�V���Q�y�e��Z�@I)2��$*�"Rݩ�*Q|�;d���z�4����K�ڟ�:��쭻��:ش5�E7���br��
�l�h
�|��i4�|�ht��Q�3y^E�I��
@���6�-ާɏ<[�܍>��1�A%��{l)���:x�kf�dz��ere������3��+2�k��N就�i��e���wz���]�-�V,��^g�RQ�Yq8QrK�i�ē�sR�t$K�IIn�M����9�nA�Q�����@�$bm�X����01^K�[x�|��}�(�eL�iW�G;�u%啩h���D1��!�ϩ"}�E '��f���*㞔>�Т���f6��J�>�|��/V%�!},�>n�b(���毗9�&Q��\��^l����˝4��&M�$�]N:9*Q�4Gz}	f��c�&�Y��6Q���,�rv�l��^h��8K9B]�S1��9k%�.�06�D�v ��1&�J�����q�Q�k+��b9|���:)�s(�c:���#�a�B���
�\��%��:�`���*Q��L�����ؗ�8�~�zn.�%k~�Rj�~l������Qw�O']6M�9�riK���o>���@�{����/ց�T�#���x�)�Q{�&�(���|�^W �e�6��uX�e/�)+WGY`N�J;�BvA�Ɣm�m� �����׈���V+v������t�ݑ{�ڭe:0AdCL������j�Xm��������sU����d<��78�?<��k�1@�nx� U�C̦�Ȓ7I��D�h��^�?[!�t���3#w�],F����KmӀ;8��4Q�ڧ8d�ӈҠ?l�A�]Ԭ��K9��o!ֻD�J5\��lT~F���!���wؔL���.����o0��i��S�G�y�nZ���l�Z�x��٠&_�_:L7rr
Sl�ҩ������50[3��-3	�a��7v�XU��4;���&׉��n�/�Z���T����h��:���le HGқ��PCp���w����7�h�(��r�M\�5��� J�S�:�P���y�<WT%�ˠ(a�ܽ�����X��#6�<s'�U�����ܩֆ��<`�>�GM�Z
TV��k�9��X��@]^0$�dQQ��x���E�?��lg�o��5/r%e�� �����|�蕄��!h����4���127�!�V�c��$8���_�-jrUIݬ�b�,q|Q�Ϭ3/���:� q`�~D��i �u�7��*���}܆�Z��d�Ą��;�Y�At�~������g���?$CΜ�����'�[B?��d=/zl����j�F�R/K02 4ͣ�|[�;"�SMo���iIJ�K�{�I�=w#��/"DX�iֹH���!/f�.J�M���A&CQ_���+��^-s-��e|�խ�=7,c�ɂq+'B߈9ŅՏy��1��H��mvR4�6V���'��|�&(�B1����e	i����c���;��%ӣ�'dF�j���2�DL�!ۦ�e�7�-�m�I;+'~���&��'8Xv5P��:�q�Y���+�Eb��E�����p5\vN��Lw&A�����L���v�$z-�[��{w��?
�T.���Ĭ!�o-�a��7�;-R&�[�r�:j�����a�-��t��������,��R�c��PK   ��:X��yD  4E  /   images/68f8dc93-d533-48f6-a1fe-8db98063bd4b.jpg��eX�Q�-�-���Z� �����wM�R�H�Eŋww��	��B8����}����ޙ�O�w٘k���\3yXxX<SWVS����>~ K E ��'��G�x|0q01100q���p�q���p��I���=�xFLJFNN�ODIEAFEBFN��4��:�O11�������N 1�Ћ��xB��N���  h�h�1�ړ�1ba�<��{,P���	��Q?�z|� �$a��"}��ٍL($!�E���\g�U��=�).%5;�s.�b���/��UT��u����M��6�v��=<��}|���>�����NL�����=-�G^~AaQq���ں��Ʀ��޾��������s�7`�[�wv���g��W׈���� �h���q?�z���������10��H��`�s#e
�!SHȭ�z�"�sJn�>�K�*����?������쿁��E >:���@�;x�|	�E>�%���� ��+n	mz���B�� �'�a�+IA/���< �R=9��uY ���L|bm��g���?o�͂���9��6n�K�}�{ޤ+���I��M�ߚȷ���w���ЏA��L�����;d�n��$��=��C����z�Eʅ��
�j\�^.V�F��w�� �=��/� *�HV<��{�4�5��d�'�D�b�\�x�3�v�/��v|��Lp1�k� {�G[����p�e��:rW�����l�G���)\��\{Iq���<Adv�:�}��Ah0��y���L� ����U�*���ь�=�ػa�=��u��MJMou#Џ��B��5����]幔Pt�o��Vg� ψ��L�rg"bz��cl����:����/�#��!кU� W�G�����=��m�f��m� ���/	Xj�ۑC�%��nr��4i�k��`�Ҋ?�(����Ϗ�wb����k���w�Դ0�/yNx�+^�$'�a�+x�`���`E��gq4_���C4��V�U��&P��?}��G@�q,ɋ��J0���
�Xo3���U1�ūr��"���gU�n�o��U
%'���X�m��SAy8a���Y���/�'K��(�wG��9��6�y�����V|�o���]�A!�)�6����T|��l��
��3n'�mwF�k߇\�r�ty��o��Y��Pt��r�L���7U�) �EGa�5�M?U	�<�*�;~���ذ�����6} اm�b}+�A�N�%)pE�?��yQ/M��}�Gor����s�+��"���.X�cA���l��FζC���D!�JS8�vc.[�9D��Z]�ܟc�U�b3�~��{��C*$83�֓)�FN�^&��;��L�(<?*�M8ý�kr�f��{V4z��/z#A9�ͭ�~�Т�	�4�W��\�^�ӈ�"��\�!D��l���}��i���P�@�Ǝ���'���7��ԮZn&�"����Nbz�v��0=]U�B��,�᥽�@E�9�ɤI��������h��D����<�^Q��X}�����2��7J��k�����S��l����J�N��Y�C/����uK��<{w��@뎔��K� G�� R����i�q�ِ4f��#�%���"H�xz���ŜgUު��>6	�d��0bβ�$r�#�rP)���7�ʀ�?]q�i|3iI�����BFkuU��jT>��(�� q!�:�L�[r��vN���fxP[���U�]0�h�1�c��E�ˈ���C���w&�`<�o �Z�&�j�D�Xhwތ3&S�P�^��n}8�p;����nʯdR����I��X�ިK�9P������A*ω�M��{/U�qal4^�
�:��z;ub�wR������#��*�@_oz���D%����Л*1Ff�����;���j?�em=�4��>������Q���v�����{�#E����w�+Ko1���-�W]�}
�09]�D��K��5O�7�5�SQs�컡�f-�N�?�R��c�"���H�5hR��-_)���;QԾ��i~6Y4��{�r�7�I���O
OC7+#n9z��kۼ����3&�M0neL@l&b���s1�=�
�J�}�k���>LHp\�A�1\�a�.�<�U��seE���Yst�K �/��L:y�i���1�Aw$tzEU�^��ugv^��>Y{d�KC__%��j�'I�kGB|_xn�N�x\�0��o��T\H��3����o�ԩ�b��{d�&:�������/�h�ca�N�����Plh�v�]�r@�1nM&�.��6�%��t����^���V��7�m��}��w��H5��7�ϳ�R�_�J�m�'��;�S�Vg��Mt�K����Oz�u[�|�����8M�D�D�7��$�a)sx;���;[FZ��"�e���-�CITx殇��%�����>��
䂌ܲ�u7���잣5U���/�Z��;]���2�/������[���$���b�]���
�8Hu9<��0Kj3��i��Ø}9�;ݪV����9M�_�Lcqa6[/Y�<T�G;��fuN��tN����YB+�������*�l�=�������?[�;�{����/N׺V@�pT~:4zS��"�ܱ�������.i@_+�'�e-V6��+_�-,-!��G0�(i}6~%�*X��2�Ȳ'�9P�������dW�d?q����D	W�xU�'CnU�� �����_}�.��vr���+s�G �p�	����4:��ۅ��W�6�٨�H[�B�2�==�����T�e�@�k¾C����v�����D,�L��KK
RtQQ�\�;#�3H��� (p��v=X�j.�C�U��'�PZ�2~�N���bM���x�f� Қ��r����T1�?#j:(�5��Ƅ`ҎM�I=�=�*ç�W/_ا�W�t(G�)37�9��)iگ6�Z�����;UsG��`O���;�4A'\���w+ٍ�6pO1JI�ә����~!?��
I��r4�?XEs< ��>�T���>��}v��-*$��>��p�BQ�> "a|5���x��h��i/j��q������EaE����HR�9��f?��O���/�%������ΐf��
p)��?9y���B>��F��E
�E���\j��c�;�}�ɰ�=�\^#߂�JS�]z!�HA��#�;�i��-kb�������A��/�x���Z�f(��>�1��������!R<�@~���z<�}�Q}RFh�.� �d�i�e�&*��?I��!���MA$t�p�~6ٷ�1�-���=�,�_�yz��@����8i�O�3�65����Ԣ��du�]�@��_�v�R$d��qO|�����!���f���/&��G�Ӭѳ�s���M�iT8�X ���u����^%��+��hSM��]C����;W�̝	�o���5�(��C�R�UVY���!1@�������'�}����j�h�Y]0WG�v�iV!4��t����2e���Y*C#A��fLX�Q���"��r�O�V>:�j5��~Ά�m&�Vq}�;Kl������A��������1�l�7�z�Oڍ�������iռɷ�*[ꁽ��b�t!�7ҷb�|;\ǟT��J(LmY)h�[����"}6 �f*EjoߵɭzX7.�<�
"�k�T,�^��ԡ��H���x�2Y�QUb�G��"j�P�N�/%9�FO��}L:�����u�za,�:�k�4h��܇{�>HV�q�W[a�T��o���.\�%^��^��R��=��Y���o_C
<1GcƵ`����ߐ�G���J�UR��$��ך�����N��.��Z:@��H+$�Oe�Η�`S�>%�C�8�☂q�-��R|�T��tp��nv��k�/�O���F�l��e:&I 1BY���u�S~7�"o��B)~(�J�X��eF�����WY�}��5�������K�]��v���0�倱���*`tM���Pw-BeH��N�����8뽋5���9c���c[&#��j�Q��ڶͲwQ���cî���5��mgh��@Ja���ܡ<�`mq��r�����mv��C�U����|z֖���;��4��s�u|��e��!<5Ѭ՘"�u�T�N��b�X�c�D=Ez.~�?�j����/��G4F��#�Y�sQ�4;/�Y'��F��9�R��<�Ϥu�=]U0��ȓ�6	�4~�{���jjfc��(SP��.s�*ꁠ=�1n0о�d�����q�KF���q����i��@�ǵ�i���5j�a��u��2�+#�+b��/F_���H���B������
���ͫ>>)�`��ĸ�,�(C�	=C]����#m��M����v(��;���2	 ��9-���!>������'.u�/�a�O�I������*����7P�l_�ޢ�aO�S"b�`�VR�t-�y4�XU����M�a]Z��W����� =�$����_4�H�� ��=s�6g/�Kq���Vޥ+�<�����Ƃ6\>���}71-�������f�=�ZA�!�6�f�&=�e�tܯS_�Eq�Hg�!��<�,Hg�'
��G|���h���y�ƛ�l�s��4%�����������5�����%�*sBbo�$oin�,k�g�U�)��$��ָx¥C���-�wei��96���f�.̙1��3�g��1�_�n? ��2����L~�;������%{>8�S�-А��h�u��P��~���Ex�`�X���� �㒒��sè�`�WD��ԝ9����c���|k<���1�4������C�8XP����4�[��
�(ߙ�=�N��Ԅ���xv��:�ʪ�)���3�٪HǙ.�,..r1�/�a�*�|�i���oy����U89/��0p� h���;ϼ��*}  'P'�Y��'����@����{�o̥!n�ɜΠ_����(��Eh�T����H)N�'G)Tf��p�*7V���꧌��$Z�^�.�+t{ xҼ�A:�׽4��>@�>K}o�,AuK��������g[gt��� Q��$������&x����k5&�WdPV��b\��M���EG���=���Ny�@���e�=�[�~��l~h��n�6�Mi6��hN�4����-�GQ!=���Gf����ҡ_��V���$��}Y�	�17�;CV��q�?�T-羚{�O.�u�%�j�=�A��P�i1�N�0�3R��nq��Ӗ��n��kǜ���|��;5"�B$�%u�%���1+F2ǂm<%���N-H���p1<���ӎeB�DױĄ�#ȉp'��}��β��P���� i�Er�"c�BS��	8Ve8��e �uY6��*BvT�Ӛo��$��3�c���$-��Ĳ���,j�$�#�5�5���۲Z�1D~'sU�����U���|��>e=���2K$�B�>��(��H�T�x珗��ϖ%�I������h	��6,��J*��"eG�c��e�fUr4���Bd!LJR��R!�~9U�<X�to�7o�H���־�/�k����i�Fo��dɨ���L�i;���!)E��^���N�`��68^�CP�\w�0�1��_�2cbl�G��8"z���=w&!�W57o�	5�F!�<y��
N:��!��FLG��t�Zb�ü%|�/} I����v�p� <!���2]#_[P���d����`�;:H����t�c���'�X�����YϬ^�i�L��7{u�¶q�u�غ�HKB��x��$)��NV�kK�-���ƉxJ�T������`�ǘ�tAA͞���F_�Xz�0����cL.�a�W�M]�}6�;b_��,�{,;�Dļӵ�2V_�H?g2�+�!
�8I��vD?����l+Z|F�k��r�/	�n���y�o*~�>/lRf�t7�����_�T]�N�o�(�� -l'&9�� Xj�n_CȤ�E
�����~$�؀�m��Ia��J��?��'	p����7���x�����(��Z��6���� ���㱮?W�3C�UE����;��Z�	�fD�&祆Vʯ�"�G�w�웹oP�V�m1��z�]�] ��;:�KTh�"���V�aQwz��-��+Oi>��r2uNV�)�݊��P��ke�M)�b���]T����dJ��##���􇌑jp��
�@u�f��X��F�-W�Y_��|<�w��_5V�FϋJn���v��V�S}�yX�~��>�	�D�ux��"��[4�Һpn㩓i<[�X�����7��pEc����"�7��d7&��3@¹i�te?eukN{�L�%i�0�S��;�_��$��s�0�p,�^w���9����X�a�5#��Jk��ؖ�6A���Ó���,m��q=�	�5�;B�r;%��VM�ܼP�y��]\������ @��u�y����4}j�`^�[��u�w?�>K�n��"�E>} 0
? �Mop��{�i �5Z�,���}_["Ѷ��r�����3v$/C�}���Z�	yѳ�����Ӣ(���GGƯ�p8Fb���������7��20�
�w��̋W�
vb�����(Fڨش=ؓ�'�U��b�ܴ�&�u%�Jp�Ia���Nю\\���Cv�˃�#�-���Un� �u�#>������.6�o<�d�U�Y�jQ�\;ܦ�(B�;���9v�����<�3	!�K�*�?8��E̼������i+G��ϭz90��#�\�!G��=���ML�[�L���j�n^V&����j��YU��l�E�j�H__��B#���nb�6�+Z�m��>���t���H���t,���j�s8��Y0����P����%Ȏ/s@1M�1�ft���j����o�ܮF�ov!����$7��i͉� ćP<�3q��ݫ)�� �����2��MsY����|����/s�»>~��k�@�\G���j��y/O���-�f@YTUc�3�'5F��/�5z{��h��9��y��U";�D������߁9������,8+�~�H��Q!Ѯx��G)=�|����,}8�^���{5�j�����x*��h���? �H�F�
���/�S� �Pѩ�[�RI��Qݨg���c.��fE8�q�VK�Z8�G����[8�&(L>iT.��������ǿ���k��o��hS�1��)l�pQ���	��y2�,�q6�~Ԗ��
�(��2�Y�tHDlN�d�#����t��J�����������%��6uńET���/����ۏv:ԏ.��6Y!Bd1v9�:���۩F����[Þ�t���Yh�eQ�]?�x�����^mͿ`��W�A\6rJ�˥��ӏ��>���:&~S�dy���:~���7|l�S͢�H�\��DW����)Q� *ˑƸU����M�����	b�l��� ��T0�
k����ī�Y;��|����u��� g��G��S"Y���0�2ן��{B!GK�ђ:�@M|2kBu��Bh�͘?f�Ja�R��S�p����*ϬZT����[���G���c��5�;-RLb�<�˛�.e0=Up���rF/P�.ѩ�>,s�f �.S�������:�[�	��Qd�m{�˵*{�3=3z{ܬ�D!S�ѪI��1��W1 _� ��p��xi�\����N�ł��&P�����?�"��(2�O��/�Cr���~0W��m��l�iI���K��(�r�i�4�Iũ������{Wb�e-)��k	!�%��J���@Q= Ro��	0���E���;qd=�F�����[�z�@�~�Ӭi��0��v^���ıإLT#h[_<"uz�_�6.I����祄]Օ�_�2�����)�(��.�����DQ< �y=�VX���������< ���U�
�=LY�6��8%�v�dI�����H����(7//�T~oy���gظ�����b�c�����b���gOy�(�>�h�"sv��[��@Rϓ/�a�&z�K
g"��=�L];�mv�X����zGE/
7�J�⭄=�9��� ��{h�O����%�R���f�nV	��\e�
L_Tڝ�G����5Hk�hG[�����C��f����v	��ĀG����R��w�8hR!M�їWxG�0tѕ�}z0������ڛ����K�W2}߫��/�<n+��]�tC����A��u�!
�_�3=稚ͺ�߷5�z2U���gpũ$<,�m&�_	Pj�w9>b���ᖛ�D7�d�囻�v[��<�"�PV���#\2��uï����ҠSE˩��;ӑH��S�kr�Z�z#����=j
&V���j�Mj!"��x����U���}�/������=} T���O{�ʌ���?>���T�l<��p�ߪ���9��ۀ,Z����7�HS����<��Q�N��.�,�`2V�D�ש�G�
��Z����t؝�?���G�=��۞0�yK�(��tb�C�4�gH�ӌ]�O�&K-e��pH��&?�r$
�D��7�C�ךs@�����邧n�[�/#�6&�ޟ��|�b!��ۊE��%+=��ޣtqH{�Qh��I?-�=���P��5=�S۵���֖��}ԗ�{<�;xT�1�IOi<�_�d5㮲�&�j$h@0i�E7���'�U:oŢ/�5��bj]W��0��Su���OD[��D!z��.G�l���h�m	=��j��c�Iw0pc>|(Mt ���J��x�����V��%�� D�
�?�oʗoq�	�E� �>�O�/�u��׭���ՉV8��y��Y�d�u�hc4�?��%P��<�+l�h�l�H��K�K^�����O�"�� a��U>�sǫf���~�4#b��
�xR҃6M�gL\B�=�~W%�F4�"��Ț����e��|�
M��We��Y�h�<�1��b�?Hٔ��]U۹�a��nY�h�ND�$�Z�E��t����@'���O~~V��ç��.߰nѥ�b/�T�V�ž�cH&��TR��7��8[�H,�ۗP��IiP!�R-��4O��!3���S>��S�u���<���c��Q�]���i5�t	k���|f̜P���K��#�B��Is:��U��/�K��a�]@��n��K�(����!�!��d��/�y�?D���J�� �>�)�����VԿl����^Fym[�L�*��M{_��R����C�ʩw����'qKr�:���}+g6��N�{�����~vm����6�JL�Z��ϯSYS&ѥ2d����� �; �[C�a�Be�M`�S��q��5�Y�����ͻ(���p�|;=¥�$+��!���J;�|����I1�_�0=�I��m��A�;����J�oi��:�0֋��옼���Jj8�]��o�p�Pi���.UO+cX����7R��f�h>i%�x�ŋ�Ȣ�z�'9���'�Y������;0hg���D��f<��@�^u	��+�����ª�CZ�J�,mۖڗj(�'���1�y?�*�-"G�P�j&�X;tXK�<����b[���EV��"�[��J4���� x��}@� 0&�P�Ǒq} �@" ςY�e� �Nz��K޹�.�Se�}�j�៮DM�
�-CZ�_�߃�b��y�f3R:����&����I:f��/r�+&�5�����A12�Y#@|1��[4�bD��&�1��n99ᓿ &����20��z��-����[����ßd�>_X���~{&f��tF�å:׈��'� �ƫ�S+~�+�N7���c��ؓ����;<�6��-|T�Ʊt%]��N�6^Ob�"HQrv��32]i�q�O�禙w�����3�:�Y�*�o�0�ڿ�HbE�Ʌ��\8*����
 �c�������}��G�ܩ���]�\�?��1�C�Qp�g���i��D�kM��_�q+�o����ar����W���1bô�1�6ӝ� ���w@m�e�h��)��t�W[#�//xϣ3�-�r��I��;��,�#��<=:%,*D��׎)Ø���b;޺K�5Q�E��%�%�:v��\>K���/bw.:�O�
4֥�R�$�y�'�||H
����yV!Z�P+�?��X��M��;|x����������i^i����nM��7rg��#��C:n	�6h}K�\�-����Nh`83z���G#��B�O�׿��B<8��*y�r�.�b*���[VŢLxf��EpO;��Zd -�c�\�v7��e�<m�|Q!��"��GV�s�$u1~�~	5���g絡�n��-��6����4>%�����H����Ck�#6���n�������\����٠Kǋ�w�g�J���^�⭎"l� �e^�r<K�g���]�#(�֯�w���ͷ��V���*�m���f��|�˗Ջ��F�M~A0υ�1��w�^W�|[/e}�C�И�9<w���QZ���G����o�wU6[Y���(F��i]�8�B$�Y08y��N�b�U%���nlaB��b6B����P�QQ^���z�±����nM���[�zl����K�{S_�O�Ն���Z!W�����[�HȆ0\n��M����W���;��L���%z2V���s��K��������곜�p���KZ:6K�9f�Uh�p��V�@���.G�o@#<�I�K�G1l�.b����6G0u(9*��c;�P�HyD�F��SD�.E=�M��c?`���-vKN��}WCp��z��k!���8���ϣ[����2����D#��v�^ċ6�z��%�즽�t��^��e�F�N������f�|�8��{���亝^�%K����W�ɽ��4'�I�O.��eNdf���Z�!R��I*�*��`����i�N�#(r���=y19*]�*�c��)�9ݦ�Wk�>g�O��c^��Ǆ�Ot`䙴��ICExٟ}���O&�[#��C���UΙ@���>�&�/��X��_��fq�#��}-�+
*i䛃�&���?uD��>Y�&���+�7ơp�n�f�Bk�<��E��
I�Cv�SRk�;��طsN!�6�������sQ'��~KwJ�a�#	=b˳�X�~ �����J8��=��Ý�9��L�ہ�Dw� �ّ�$Y��$�I��Xn�p'�gLό�< �R)��!���������ڜU�c�"m��Z�l	5�l7r�vT�q����p�� � V�]���O�z�XܻNR0��u * n��0�3�(���~�;I}���{v�c��^��A�w��yTr!�O|�,s��w/|u�b��̵K��<��y0b��:������8����#Oԑ��!�(���[r����?�c2���߹�Ig[+����CW~�Uo��/~3�h
��Q����#7��%m�]?��;��mK9a[j��$��s,N~ţ�U0�U/Ƌj�|J������� ��3�CE1�z��B"�$��-�s��������<z-�w��8)mZ��l��ߘ;��`���*�mLW�5�����sY3W;��+��#���p�km��@�k�ct�*�γH���=ѥ�i����/�|�>�h��+�L��1*?�ʊ� 
�v���.2���e��XR�ja?�V�X�2��^$�A6�lg�5����K��/'J��K�o:�t���iV.$�2}�]��d��wpK}�I<�YKo�sgQ�q�����7���$8ᣄh<��/+�k~��m�h�@oT�����_YǗw���7юJ	���\���6~���#�	�i��ً��ޔ���f	��9�&�T�*�<�H��Y�4{��Wѭ�͟2q�����h .���vZV:.R.��;O\3�Uee��(��!�Nw*��s|u)-�v�����}]�6��(�~32�Æ����`-˄AL�	x��?W4��[\5�/<y�U���耀���y���u����<:����Fojuԟ�\�颟+;�����ڊ"������/�}�4�F�N;��7�-��8��GF\�j ?����.��7_/uE{E�>!H�U��#�� �T��/��;��������7��>>���l�}8!4q<P��́c�$`����3��Z̖��e����(�2�y�Nq��w��B�w����	a��0ޱ���$6����ojџ:���[jү��H�S�~Y�׉���� �-~�RC �a��k4�����;��QŎ��%�ڬ0ܝj\Eδ�;�oGa&�.?�4���i%�|7�	w���ē��(�O,�;�QܖG��v�bcס�4=2
�2���ۏGw�с�{3�=�`�%a/w��&�L��Yv �B�.��9��w�-y��)Yi�ǯ�^���r~�E�3��jDǺ��<��ͪ�ȅ�����W�%T�������o.˖�΁� .?���	!B	"EZf�.�����t�"/����{�:�^3:�qI0�/��'Ʉ�7̉r�,�L�b�4��j	���e���v���RE�'k�Lڪ�j�n��� ��3�##�咎_|�䦒u�Ы$X
�������G�<���vZ����T��9�yn�h�T������)��8p�E��z���*���4���@Ĝ�΀l#��f{N�^�n�ˆ9e{�vk�W����Bŗf�%��:�g�L'Ɖ��k*V.����V���oȂ�k�5�/T�#�"���+B��-)�^��!Hw3�i��*L<���G��y�u E�C�^�eHol�?������^�M�tu�� w�{��O/�̆���c7t�oף�zn1[�W�L��d-��κ����7���8�jI<Wo�=V������,!=�Ỉ���5������P'�3v�����Ybo��㥹 8kѼ�P%���oU=�"m�El�v�i3H7AQu���DI#p��Q�R|6��.~�Uzd�ʵNNٺ���	:�y����rf>�R)���IqD�� �c��V�6�zL�="	 
��;�1[���2ߍ�:=�Vr�c�y |.2��q_�3�Yk�o*��,�֯��fU�q���Q�3�s����5jbduB�_^6K���婱����6�=so�cS�����s[�8y���z����Χ��s�E��MJi�	�=\;����BK�^�V)���쬶ݧ\,����_�q��y8���8,'�/(g����ѫ��(���F�vMw�z�O!�,E���C
��T9��-��Q��suM�ص�%S�� .K�׹�>R;�C�I�v��X��X5}(_�0�����jgs���֏�Y��+�1�������]n�#F:~�ab?/���	v�Y�q���)Q���v���_L>���d�u�M|V;βo̻$���8���X�<��~��ݮi�D�Fro�d�v�������di95��UNe�R�p��*�^��p�	�~S�13l@��B_�����O�e/�/��X������2L����M�4�X� n�_?p29W���@�z�w�͵^<N�-1�b2�D�k4ڌ�e���Z�/&`�볆6U�؄oę\��4_!�j����ę�W� ����h��v��j�.X�d\H�GJP��-��Kcx��ۋs��y�B���ǐ�/�6c�BBb>�̷g�E0O��PE|�K��JoO+���}��>�y{t�һ5^9ր����ɬ���D�ޞRƿ�o�J2/>eZڜ��/6�m��%R$��$5޽�^���i9b냯vv.�s)q������q��,�7`��S���D�}e�,��&� ��D�(�J��.T����m�'�k3>rj?�g��7y�2�>���W�A̨*r��m*��9�n- j�xQ�>��.�yS�$�gG�K��\ݣ�o3��oO��Q �	��$����i���h|����?��|�pg8!�9}Ly��&j��b����4vd�ȻP}�X{��n
xcD]��,~2Qh��X��,��0�8]���ƫ���(u�E��̃��M+�7~�W,��Z<j�,�@�b�f?��.5�4���]£��HQq���`a�R�7���ip�S�o�G`
���C��]��:�e<����+�F�1&���8wxVB�a�k�A&��ld�5^��v��y|F�2.c��nBz@-����+�_}��xQh��7�C�#�>�4���[ڨ���~bdSU+΢S3�#A�{��uS�w�x�E[5QzG'�oQ�k���S"��r=��r�����T%��w:�> ��dF�4&�|:�*|w�ye�g��Ή��L泓Ht��c��d,իMiⵏ�����{ T��m7@�����)ޖ>�l>,'�J��DE��ܔJ��XX��1�-F����)_d�8���'y��Q�xd������c�w�u�x��w���ͯ�9��uc�p�n�}~,����v�f9�lID����Ae�iޥ��?I|��I��CDr��Q�aѴ����.彀�T)��Sm�ҽ�&�Gz�j�n�D�����/�\V k�f�K�2�bX�s�u��Zy���ĥA����S��7�,�3�x�U Z�]B=�.eL6x��-���ۍ�0(@:r}��H<D@��[���5\j��$����M1��r���g���Б��ק������������f&Z�̒�Kt����n�T��ƒ9�'=��*o���8�5v8�Fb������(�	O.���%�ǋ�!�a��Y}�1�D���M�Eʄ�|u���&���5���J�� �� ����jb(g�TM��*���N���Z\dx�}a��fUc�P����P�BTmȨ�u�V,*���y$=@'�ؙ��L>��.c"�$�����޿H����y��2]/q2t2��(J��ո�D�y��mR@x�#��Q�U(�v�ł�t+���d)�L^T��ҋ�)J<C��9�,�:��MKM}������K;��F�d}��=�$6��z�������t`�mdˋ�bR�[(�L��.���!�݋]%Ca����2�$���׸j���>=oٞ [��e�t�j�������S��E��BT�
�Ah���&>��H{ݞ{�h�T^?ݼ�rۋ޽�ۭmQ+�
��Oڏ��5˾z����+j��v�"Y�9�}��y^��46,���o�T��E����s| ��b����9P6`R�2bRS�r'�� _�E�~�r��ɦ�;򲭆0�zK���b0�$̯fm��;/�D��o�e����?��dh�x3wE��.K4D���|���F��Ϭ�qj��P�]���I9����vJ۷F&ˈ�|3�4~j+��j��qa�e��٦�]�>Su�b���qU?�z~:�Mݤ̻�o�= ��*{ר��֡���&�3�	���F���cIY�$�����df�� (߅����ڠXy���ؘ��~w��49��u/%�1u�d��Sn�C�	d��
)M��S���?Mb���;Ή>2�y�ӷ���z~�B�5�B���ٳ�}	q*:Â�ޛz���7�i�	}�[M���Q�=(~���P��*'�-��B�Wk9�a �Ħ�����S��U������:��Iףjd C�W|q�]��:��/OU���ʯ|-
JxqmA�2Y�Ү��u5W�3��`Fԏ��?�W�3����'7�*?��jN�E�x��*p^�������,�T��řݩ��Q��akx�=Y�:p|���A2���~�#�r��:�?�g���Ҫv� دЅ^o��\/�"�8�� y�`;l�T���X�;�W�p��M��  ���<���H����]t3�S��&�
�͵#A�S�;�;��ҥ����72 0�N:6��5v[���/Sy`���R%��}���!���;I��l���W�('��-#׻,Ԋ��Xpfn��m�T�jnZ0��%��0���Gj�� �~��=�Y�Yf8E����_�_�C�a}����nTX�_$y�.�c���1	ː�dh����k�$����ػ�&VS�*"�#QF&ʲf�0V����>���N���>�hg�k�P�MtZ2|���5��PH6�oe�c���kRޖO���VB��CT&�O��Rd�+i�[XX�Y�>J��@k*?y�qG*;�m�i�P���8������D�K/����3�� G���3��V�;m�Ł��`*����$f^y<Z���
��؁6���:��=�����Yh�E�{k��]m I��܀�4ۖE��]{h���W (���~TOEt��>�?�4t=cy�����r��::���+���� h};������.�۝U�<��F��l�6�FEh|w����6�5�߬L�a����-�"�rz����>���CL�Ɓ�iZr�fm�rř��,��f�O�߳���+x�I��GĿ��,�[�C�)aֺ� �~<�����D�n�g>�m���-n�]1^��*H=��2���Q�|�Ƈ�jޫ��Ym�)PW�89l�B�
 �Y�|�	� T�� `}9��[��)BYx!�� ����E@��XQ�RJ�|���(��<ʺ)����Q@|�)x�4zP�(>�úe��ڪX[>����H�Ȁ�V�@�U١K��J7�w�t���=h��������N����L�eđĪ�V e�v���떍ky
�
H+)��b8����i�� �[Xl,`��������c�(�f�j^����k��>����I�²(aѰA�z֘���� >I�i����1Y��t�7W�T����.��D�T`����δ})�� ������(�>� �t9�A�ߍ�3o<5�jZ����m{4tB��T��A���Ydk���c�=�ڗ&�3��M�u)�kq��6����}�8��{ջ�x�1ț����֞I�؞�OG��<=�-2���ݜ��DJ�cd�́�穨�����B�.a<�C+���1�M�߭ *�p��m�A
��T*"���Vuǆ���Z�R���ak�U�7��G�V���\c� |�4�Y�sɦR�w�~� �� ����xG�<��n�P��PK   �:X��S�  �  /   images/a8eccc96-6934-432b-b3c1-5526b5feafa7.jpg�WgTS۶�!��.D�*Ҏ %"��  �(��((ңB@i��A@"M�J��H�5AjB�ϸ���Ƹ����k��k��׷�1�9'u�:p_506 @ p�� �	@ ���4��fzzV&&FfvVvv6V66N^nNN66n~n�>>>v.A~� /���# 0m=����6j��D�`�i���Q� ( �@����������F[P�Ё�`:z��S�f�i� =���.�	��L��C��$0K\�h��G�Tq����/ ($,%-#{欪��5.�]�7042�jiemckg�����������a࣠���(dt̳��)/S��32�^�y[����}IeUuͧں���ֶvl�7�������ѱq�����ϥ�_+ĭ�ݽ}���o\  ���[\<4\t��`z�߸@t�~/�gWb�յ`�}��i�'̐�I�,*�	|��}����x)�oh!��{��B�/`��� y` +��	��V����Ջ\�!h��> Դ���snaF�d��Z��> ���ć�@L�|C�s�8m�k�H��v��bƞEr(�ߜ ��<-j����m��P��~* �VD3�?�i~�Q3��C�:��P����Ʀ���S�T�_T�`����{�f�^DT�I�P�=NEX�k���VT�O��5a�p2\̗��^04c�N']�їKGj}+7xx�s��1�^�{�0���\S �	bq�᷻y�	�*`�P�R��h��Ǧ���>��?�@��z�k2KE����W��	b�R���V�)yE�L2����u�&��^�t��\+$��9�������,�J>EZ$�1'!�o6�����?��Rt��ߘ2���+B:�'�`<_t�������+sL%��)����Ñ����%�w*�|}������NJ^��;�^�3���j�P�t��D�kQ�8�?��6�ɜ�l"]�wG��N�\�R"B�(/7��8�}����N��t��9���rY��S}{����;��^a*��;g:��e�6��~㊡�1�t!v�gWt��
m&`�"��LT����|s�D�Q:e�}��Zw;���(:V�O��"��!Q��?����������U�+�A��t%-�4'�?e^aF/��,�9�@�ZQ&m�tjn��ø^���$���������4m��@�MCZX��!� ����0ţ���ו��|#,/	Z���Z�|1uX�����q�C�Cs��fܳu��\������W3��26D2��Ӫ�4�,ZV��A�XOFvZR�c��|�H�KO�Xf_|���OD��xm��V��b�t��}	�I��U�-�)
y�ܟRr20����p'�cez�a�+?DtU���D����FBհ#Z��pT�y���Gu��o_J��>m��
�G\��4ݞv�y�:%�	�$���Q1fUr_:yC}�Xw�E�ڛ�N���r��߱���|*�u�.l����/S%C�����|oM*�<yu�\�~\^�n]Y3(޸2}�	�O.=�ݗY�D�@�v�Y�������^*��!H�zf�����w���eR�hS���!z���x����F�c�Eh<%ĲZHA|��ku����Wb"��ND3��|;5�;S������b�@�A^��\��|
�
P0.�˰$.�q�E�����#�v�Y���� �Txo��y�B�J7�.�����g�Ԗ�ѧ����v���\4�Mr�\H��l>�hm��k�������}��ZU�j�eO�[.��6Ev����a�3h/�x�$���2K����p��%�_b�S-a��E ��둲�ϭd����u)�Iftx�(�7�D�9�#��u4Oh�Y[ju�ݏ|܍,�� ���-�3��h�4É�Mӑ#����~�u�	X�+��������Ď1=�oT�u2>� }��Ӧ��v
Cu?�Kf�+E8{~���E0oԜ3k%��U��?�2��k�Yw7B�y� F<q��`���m��DbYԶ��z8D���֊�#����U��6��󇵤���h~)Y9��D!��>���"�e\��p�B�b!�s�f��։�<��Tz¢���S�N�?�q,ّ��� hsQ�b���6��8����-f*��D#�Uy�^�5�����Ƃ9/J�Z�mJ���U��{BF����rR��#D	��2^/�}�W�k��?��Ҍ&�Om�l�:�'���	#4�P17���*��fW�Hʒm�w�KRE:��q����D������~
Z�D�A�F�cv�ꓴZԽ�"ֺ�{��]Ri�@��p��"�_ò&嶌�����aa-��MI���]�d*p���X^2�ͽ���Ɔ�����cc��2+.k.��V���/�-��L� ���وc��Q��pZ�9�����Qz/BI'G.x���r����|�NT�F��JW����W{�cRL�~S=G��CdlL{(w�Q����
�f�k;74Q��1�81�{س�G�Y�r'Z/^���6q��=y�V��m<���fc@#0 =r���Z
���<�W�����P��U3�2�,܇a�å�V�1Bbөm��5��M��V����$0��)�5G��6u���X<-pG�b����H�}�{4J��ZK!��<:�(jaU�U�G1�uC�آ����o���O^�{�D�zc����sPJ��(15'-��|�j�Ϯu�6��베��������D�c�i	I��.�w[��w_�[u����ђX����WG��ڒܨK��+���)XZ��=��n��K}إ��Έ�eDOa��(R=N�h��4�95r]Q���.�.]�e��Z�GX{���J��bq>[p���9��'�hw�:	>��.K�0��q�|������Nyk,V2i�fჽ�כŶ8}g�%#�HK5{�<:%Iy]恻��s�+�E�I�������	���4(.C�(i'�7�/�hR���U�hA	�>c�QEfw�5�괒c���J��4+v����i����0N>&]Z&X�ַ��`��)u��q�p��y�x�}�̓��Yw��p����T�Pz�ˠ���w*��\���2A����1�G>v<i�
����LhL���W��7$O��Qp���Kٜ�<V��g'��kۄ�SC+F�yQ��<�U����w�0V�iBE��# $D�ޝ*5dݑiK9�>GWe8ۉ�A��^��Hs�ITN�Vj�hi"�0k��#EG�g��+�OGs.��B��+b ��Ќ�gu1���c�h��X����g�W�H"$�U�6'�fʹ
��Ni�B˅�zyiv��a�AZ�����O�Xv�z)~���!��*�}�]j�eT8i��9iδ���7 K<4X��,=?X���	<��e�q9
���Zro����{��a�2�{XNw�8��<� �:A���D�W�ph��>\�c���+c"��+��>����UN�a��J�Q͚����2&�X~��X�S�Ș�ٱu8�|����H�NB'�P��#<�{Z+[�5o�m�r�� �3%���^�����7�n����͇��l�4����E����CK��TNn�z�#G*@O:���M��(�D��ֹ���>	�/�a�8GL�R��W�f��1�y'Iܟ���sJ眢�~t�3��tg6�8�l]f��]����R��H*���gtm�y��0�ɾ�䚉q�Wf���]w�Y��:鯹� Y�0��������z�'Q��+��/�N�ӕ��~"�IF�;�Ѻ�#)t/��T���ற��%:���6_XqF����Q��,QK
Vԃ
�˭�Ig���yl�QO��s����W�vK�)2�t�ŰD��f�,��9	��SZ,j~�>���&s���Վ��-�#�eޚ %�ஞ!�����?�vV��Lk�^��]��.|xV��G���@x���j�L�Cy�VNq����1��W!*�g���&����Շ��.��d��&��]����	-�4i�1hSJ�eK�U��@4v�^�9|�a�8����D��zI��	�f�`[�lyG���C�\�5Z�C �����`��U����4kJBa�vܞ���렑*g�Ga����0�!���4\���_�����O���ݹH�-Іi��gTn{~O���#DJ�N��\{���0.�b��3�O��Q�yX������[��l��V�W��S{�;'��,�Y���*%G��"����Fn+7��-�:����b�O��� T��bM��
�*9��m'O��'!�i_��gë����qdA��{��˄����.j-`����v��0)_�$u�F'�YY�9�KY������(�;2<R��_*?���NPD\��g&��X�����A*�9��PK   �y&X�,J  /   images/d5a492a1-86e6-438c-8279-421a5a29733e.png @忉PNG

   IHDR  �  Z   <�Z=   sRGB ���    IDATx^��	��[Z��cU�:�=w쑡����FP�B#"���h4�E�1��k�h�QA���@FAd�Ai����z���}�3���Ǭg�{׹�����ܪ����o{����y�=��6��dV'U��ۻ����;�'���:��j?��tR5��Y�wۚ�wU�m�w��׾�����}ͦ����Ov����n�5�Mk���~��5����5��o����f���v��-&�Znw5�UM6|k��گV�������ޓuz�5�ܩZ��d����G�a���藽�^���}��և����ŋk:��n��	�����U��ƫ/<ߞ�������m�e�?����O�>�9_���u��?��?������?q������k������ο����ߟ	2�^�������7��~��Voy�;��z�w����u�lS����,��#���kvtT5���討/_��5[.(`��v�]���:]�k�Y��Ә!��ټ��i�&3�\��IM��q�ݮ
���t��sIe�w��Gⶻ�춵�lj����?LӄS���k���f���!��]�֛�V�f��ر��9�a���t>��Mki�Ÿ��ǰ���}m';��d:��1^���,�x�)�Ɏ{b:�~����l6��v���o���� �xxP�Nd�)��g;�cQ�l�~[�~�{�卮9������f�}�y�uV�u��~�gg�A�3[�2n���V���̇�xn��0�>˞��'�<f��뽅�q�	��z��5�O�����0+L"�����v�q��>cƇ�b��W�O!��'ʊ���<epg����xqQ�!Ʀ������"�݇���!(���|V���h��dd:������{��k�=w��ƺSGc<��d"��ʹ���]m����t����l�}vt|���fM�g!��N���M�p1���.���u|tT�j1��V��Afvu��Y���'���j��E���j�=jy�p<����l7������<G6���x�2�g�u�������?�Rޱ���ȸ&�c��W� c����5��j6�����܎6��.cƵ���N���|^�%�v�g�X���A�!r���r)��M����Z6?R��@�l�۴���xtx���n9\k:����Ay�,�>��~>��`t�-X��[���l6��y㵨�f�'��|\'�i��<bl�S>������-DU)W����l���2c�0ٳ��x���\��ϻ�c�>�ރ�s�p_جi�~D�]�6O��n�*�Y�s}~1������L����l4ke�N����"�m3H;����#2���)�I5�_�_���õ����t�|ū�e7���
?S��~��ͳ�f3͓����aE���}c���F�ncy��L&�q�O;<��GߋX����)s>.���3Ɨ���Q?�8��U��LI�I�-�Q|����82��S�D�	��y��-ٛu�����5�}�M��8�?�+{+��l{ɋŽ��97X{8�8{����x�4	^���G���<
���u���)+���k��g<��GYY`���BU]�M�/����b��o��ֽ�z���_�?��������vV��?�S\ ����P��ќB�,1I�+��`�&±�20e�W���u�J'N�Qx7ۚn�5�VM�p��5ݮk���|sRg�����Z�y���U���?����w��O�m���":�"���'���QM�|�{���97��~~��+b{��mT��I�������,o{6�{����b���g^�|0�l����5:^r2Ư�<�9�~8�X��vR�NV������������՛~�W�Oݬ��Z\�\7V�:�ym狚.�5��k�f��֢ն�y�MkC'G*#F�����0��G')�K2ՕL�9�Eq��B9�s8Et��i�1��� �A !Ƴɼf���}�!x�sLg�,�?O0\�܉0s>��>��k9WP�=B�k�P{������8m�����=+8�q�H.��m�O-�M=W	� s�9a�.k�k28�1\�ś}\>�ϯ�
����އg[,�\@��or����y|
��VC0�U�����=��`��k��T��)A��M[n������&�Wp)s!��u�����ն����b�[��������猣fO@%�<ۤv5��>�Q~���\@z0��fǠ�@�`���\I��r�h��1�X��
2��*�;س�Z.fut���.ԕK������/��r��F\|�ֽz�{?P�����ݓU����B!H�̑�Nk����h].P6(ڿ����m�X�A%�0���X�{�!�3��~ؽ�S�ON��d�#�7.��؁��:�)?P���y)�:"�Z0�Z`��}C�!���Ӷ��h�:��~��@@�=�g`�/���h�I@.1�c�M�V��Rz����7p�
 {`����hغ����Uc�^`���t1�ż���
x��^����*�!XG-�� :�'��DY_zZs:��0ɗ��x����^��W���n���3��u���)��]�9@�.��;�q�{� ��c݆ `�/�~��%/�v	��Yp�6o�g�������8ܢ�~)��=0b�% J�%�G�����[��/H���l @K=��3�c��]���ށ��S4�9�#��a>+m�w�nG��>7N�G�Tv� �I-�3�� PS�P�q��اjq��τg%h����ׁ��~��b6�.�>�^��/0��J�<�c������396�n�==��Vޒ��	�6����܃ �}��^�<�'2�9�#Q�k@ob.eG����t�B ٜ�_�8�H����?������+�Nڇ�?$PYr�d�z���-l��Y��k������$A��N��Hȣ�}�=�m"`~����~��N����A��?�.AG:��?R�lv��v2�;U���g}���}���ۺ�����B���5�ω<S	�9�Ӝ�6PM4;<v��U�'B�k�	Ë�h�l8$[	!>���20��d��75٬j�Y������xwݻ��z�¢~��}v��?���ҏx	Wy�	0������'HϔD���)?�����.n9gB����H��/		??�
�A��8���>����P���gPd2"��J���J�+��������ݓ��q�c�`�q�=�G`4(�e�ښ��9�き��2�۷N���}�~�W�U?�3���Û�W?x��ռNǵBv
`���/�O��. ���R]30\(�@gQY e��[��5�T0�,d�O�d��������� ***Q8퀎(aڇ�q5(�͖�;���Ł2��%��PJʎJ��\p��3���>����![ g~:��r��A�ג���c�0^�3߇�i	�K��S�H#ß�Z�h�:��hs���2���Jثk�Y̽���EH��Lu����Q�%��2@0^](��� ��LVg~��:~�t;s��Z�Φ�0n<�h;fƕ�Z�� ��3�}�'o�q2�-�dF�^���l�P������IИ�T�0�f���Y槝�cG�L0'�,��7:�r�����$sj� 䜆��L\�	�Z����?�X.�<�l�u��I��[��\O)'fBf�]d����ժf v����r� r�`��G\;�C�+���0�à��G�E>�6����ݎxId�etd��P�L8"pp.�"?./���� �	0����>�O\F�{��DiY�I醾吂Հ ��[9��/͒m˽)���q~�wɛ���w��鎚$����'Ӏ���7��`�����]���]����b��r4���N�e_��@0p�T���8v����>i�)�ӆ�=�D�h�'����y�^�nT��5�~���,D����P�80N�v��T�����S��Z��y�\$X��Q�� ��n���^W���k�U���i4��f�Z�m���/@O�5n\�~sJ�G[a��Y3Ӓ�; LCbleOh���әaEQf����e�cFL� ��N�H�G�S ��>(��FW&P�=�y�=���}͎1�@�- ����J �|c?��es$����Oh;h�aG�'dƚ)0E�`�DA���I=����)1&�G�"�F�*݀��6�+��yʄ�}M�Tڏ`��w$�i�C�#Y��u���l��J
�g <�x�Ng��r���Y�����.�_��/��z�C̢������z���&��]U���_W_��?\�f��Y����4��;A���1����N2x)��w�&T�,�f�\��*d�6O�
J#w�`t��9��jU��Y] `v�f�o?QGӻ��=T_���>�S?��^<�Q�;�܌F��}Θvt["t���T�f`���| կAQjFip�;����iih�Y������������ �����I{�����?�8�z��ΤN�ͭ/�����-;b(�l�$�Q�"�M՝{�z민�������џ~]��/jx������&`Kh�ZlkCz��S��&(�km'.�:��[��i����s����Ԝs�=�}J�3+��N��~�!�&h�B��/�έ�u����o��������Z�6B���gut|L�V�����xwp�တ�*o1��QL��@G��/*�`lӁ3�0`�h+� �Y��H	f�f���1K���A�v�	99vD�8�N����h*ad�h��.ÿ �Z���D�,'���W�㋁��X:p
,�_�
4����d�Z��y��������2N=�H������fM97�,SS�]'8HX"��/h �hѠ��x��)�q��?"�!p�3Y<�ic\L���B���^�Hr=�)3 ��ʆ1�(~_�ƖUB�u*2��EA(~&m�A�����S@��LYS��
�s9��5>�2���r�5GwpMXR �ΜH~;�#'d潎�~4y��W�sM��� �Y=^�|�{KN;�����9����v�!V�HAS�W�$'tv[M��p�����][:`]n{�3�wd����t.�^��{;"H0ɹ�x3�r%����́I⿎&U�/�3�3�r����κ���pGm��ޡ'G�q;��Id���ŏ�*��M:���̜\�1 L0�q�2v���2�,yq0��	�F2	
򾦁�f�9��4+��O��@f��|ŉ	��Y�{��`bٓ�oЍmItv�Q	f�|g���ՙ��f�S��*_��,�n(Qq\݁�LJ��}�ɺ(0�+F��V�/YI���2��]\�P�>�N$|��F��h���+򘲏c�i���? [<�����SF{����L +P���j�w�Lt3�A��kgKg\A�%Xaajʌ0�N;�h����L��0���k%:r�9��E�YxI���Kv���/��b% �^ny�\�6�����>JiW�ȢS�J]�Ŏ�,�1c��:���c�z�_����>XH�S�"��f�۟ՄT�o����W}Ϗֽ�պ���dq���\&VΘ�("�	N���zh��B�*�g_����ke��� �Mj���n]3Ԓ�ޮK�M��W~B}������|h�A+$:�%r ʜ���P��UKe��Ή���s�C��d=�S�+ٍ}��7!���Ӷ�ih�^	^�k�ߝ	�%�L��h�q�g��z˳}(��Jş����?��m,��0d��dD~�shs=dw�)�9G�=;��ۤV���}�V��~u��W�t=uo_�֠���h��b�|@I����S�Kdh1W@�D�w� 5�S��|�kT?�g*n�5��x� QN ˳��r:���.�5'e��[uzz*��G��:;;�=A?��IY~���jqxX��u�;]�	&�4(�x�)r��b"Ҵ�)���r1xg<(�G*o�y1DT��<ŧ�H 2 ���рsv�jhh�QCQӰ'�	)�6�i���bU���R��)�g(�^ỏe/5�=(C����К���J;�l�l�����n8%Z3�dC~F�� ���$���}�1q~�]+
��d�F�01�t���� ��t۾���<:��5�-�3�gʽ������Q��8g�tQ��<�灲�rXE��sɹG����>�F��������Z.��s�H��kܾ{R�����0:�-��z��q2zp)�I��
���cֳ!}=��iUN��88;�H�� �}f���'���(Yo�QL��s��ͨ(��y���ꡬ:�:f�������u�L
xp��������QV�h^3���7g�X��樯�p�(zO`��A�ؼ>vܙ��aՆ(0e2t�A��l@z��Y[)!�����)o�g�-΢���sA��h�:����8�(�]�S� uP�^���Niu(��	f�ħ���0|B%��`��FՅ|_f�zv�&�c��&���"�̠��m^d��a���T,�2�@��S9:��OȠ���Q�]ޣ�+M��9��,�ϙR9鑦���W佦gL����d�h�G�F?圌-�p�Wa:qۘ��8 ���V��s�$�B3A;@7�����h��^8$��l��Y2�-�f��9W�����O ,��1��@N�Aw�_9u��.�I�ච��e���J��C
 ��F5��r6��N e��"����+YKF��̾�X�3�c� �($J@�t�Q7� :��{�����rwV���z������zŋ�=w`��3����?�ޟ�o������u�_0�D.�M&��g=�& ��F|���
e���-�!�A�]@�E�)�ҳZ�׵��L�S���G����w��}Χ��Z�И��������I��ܭ����N�*���pCq��.�jqx$�&�G+!>��n��;�]�!�搘��h��L��~������T�������l����QnF����˯5K� ���O�  i��PӉ5\�F]t$�p�pRS#;�}u���'�;�����<���Em��"�D��(=�&j4K�����'�׈3��n���j�����4�rN��Q �Z�	@�ݶf�:^.��rQ��)��'�u���攡
���ryPG�j�_�~2��ѱ����v�:Y!]�~�$0�%���T����4�x������߽�EJ��U�u���8�-X����ݞ��ߧ�Uɰ��Q�#& ��y%�IP;*�u*��3�CdID��aӞ
Ս�[�~EƁ*�#��Y�u#�8�v�lG����v8����D4jp�_�Hr�2���nNM��ګ��M��Ǒ����>d"X��Iq�"�h�<e�;�N�O��Хi{,�Py������Z� H�xG�%�=�F�6�F�@��ܘ[ְ����)X
����b��=U6�l��3��2&�h*G�V<i�
p����~@c�������{mw�n���p��,���Piȹ�4L8K��(H'���o�fL���� �sĦIff셊K��z��yeG	¨Ƨi�X�4��5�Bip�)驦���y H���hݮ����f�*��5�3�O9�r�����L/OO%*�|r����eM�����cjQ�M5c��e��2[�g�Z�flP�O���ֿ�wdzrE�� �KZ/e����g��u���~[o��6FM�h_�1\�,l}X#ഢM��"�#_Y��-�A������{�$�6�L��ۚ��u���z�������fy�u�#�Q�S�!�c02�Aۡ����db�֥�u��a�a��e][^r}߁��91�bd�n�Ք`�9�䵵�T$ը��X��m.����]�MFe�LQ�B����Tje��17l����J刱�bN��'���:��Q`�����%���6��t?������Q���1
�ɏ5�� �U7(6�#�M��t�b�����M6P�K���:�Qc��W ~[�Ǹ^R#���� ��dĎ1�5Ѝ�oY���BK�@>��f����G��گ����?P�_+c�v`����#����u�.��nV�ٲ��i���o�P�f[s    IDAT�]A���L�e-��P�k��O@��mT�u�S��Z �;;�C��ݨ����#^�P��_�9�_��O��=z���C7�Z��֝�7��͛ur�\p��úp|����Z,��ߥ��"��l�*��՚������q�h�sNA�.dy�e<��#_{f8�����49wz��_Q���<O�ľֳ��i4�u���6g�n�+b�_�;m:;�,�"ͮ�p�P@�����z�f9jX"!����;����ۿ�'�O����b�Qg�����13��(6�i��#!y��B1R76��F	� �/d0�)
=5
Zl�ٱFw���̺'�z�²g��lN��)��݃�ES��r����V=�����7��������uk=���B�렶�e�0�墦����2��� 0蔥�]#z����=�� j=I76��:��\�t���?�v"�6r�+"�J���Ɔ>CD�״k���q`����{=�j5��N�J�SƠgD�i����C#���vx���y�ץ��1lNư��p` ��t�4��c��P��3�/��q%�c�V�֍ܬ�g�TK<h��'`����p�y�s�aX�' v�����V
����wB=K��l�d��Y��ڂ{ЛYԀ�F�fͿ@�R�Yq=�k���	�0�H(T�%�j��;)��6P�X�tڙ�%Wʁ��lr�%1-+�aL�e�Zr& �~/R��9���e@���6�M7��D�R�����vmH�mpփͰ^��?5��
�O�k%�*����7^�
���R���=�a������dhB�缣�;�g-�g3��d�9�q\�p�ϓ,%߆@?Y_9����!Pd�gt:�?A�h{��#��� 
J��iIP�I#�'��d.�#����u�*	׎(���}�of]�e�J�M��~	t�s^j)Y���:�ʁ�P��>
n� ���X��.YѾcgf-�����P�\z����C= �؈ͧ�~�֞���������Q��}�n����>���B9|��yZ~Csu�l��j?J���3G�"9JMa����E���G�6�&3�����$�+��`� �w�w��Q��,G��AN,vs\�i���
5�2�a�<�}p�[��u����2�@&�;��i�����\m�8s���͖�)���W�����tS�NLX�sxl�N"A=&��3P��k�3������|F�7�ą�A���4���շ��!��w��1b�+�k ���l���P�-�S�I/�wb�v�I�����:�ޮ=�����?R��+̘�δC���v�ݯjZ���k��_����[�V]��z�/���}J���BQc�!T�K(��'�
�AFS�nL�@V�Ut��"�j]���)N��bs�^�+�ſ��>����%�������Jҧ�~��?����a]�p�.��˗逫��!��ӂ�q�Z�9����b��b���V���~��.��>:����`�P8`�ݝoB��@�_�����ߟi�Ώ<��"ie2zav��uQ�@���脉����ŶYx��r�0�?kF���V����c�]?���w��;�X+�X�[.k2_�p�#/��Y�g(qgLt�#Q|��SԬ�N�PX�6M�2�Zdے}�i�ݦ��:�lk��[����?Z�Q��>�C�W/x쑺��Uu�3�H���;փiw�U�;��~k]�z����w��~�g�T�x��ug=�³��-�����L����4�a���=��ˤg�Z�[I��4�l�ier�Tv��N��T�z:(�ԎF>����CC��-e3�Q��t|��o�����_�k��q�γ`�P��2�i�à�Ň�_u�WN{Q��9	�TA�&��%�t�3����!c����2 �` ���� бa��Τn�GZ���tp�q�c��95�^���	9>�HH���.��I�警=c9jM-x������L����g�����h����#����f��M཯��#"���-v�=��0{i�]b�m�R���2��/�f@bߨ���*'V癈V��"C�����0��T���Шw�ͰZ�=�GPk�yL9�9   B�)�z������J����(}�g��TS.�X��3Kt�H��ߓ1�m�����@���C���?��: L4�ھF ���zk��`�<�xsV(�84��4/�JO���������� ���t��+�Mɟ�'��07o#�����ևх:��<��kb&L��\?�>�OE�u^Ӻt��D�u=�.�篙��z�خ0a�\�U�|1\g3�	��rFf>���U��򏮏y�#<*���z��Zۚ����<)�^� )m�C ���W�F:h+=ɞ��|;��lfwq�qj��	&p�g�u�*)н[@��tW`�`m�t��Wh����z�	�o��(���3�f��I���Wwj�;+%�'�%  ye���}a�L�e�l���t��m�ܧ]���;�mZ��mm�TR�&RbUM�2�q��f��Um[`:E�<��Ur����|/������u�1;�6T0��x<�SL�_�u� ��_�7�-���r� m',��e��
zb���vU����&����+^p�����n�ݟմnT�������������5���j�(P�I����N@���!PE�i��~j���ވ#c�E�B�@{XojvvV�5=�`���֟�#��>��/�+��j�D����ީ�>�Dݾu�Y���u��պx�J^� mi�G�'��-޵rL���b�,P���s?4b��s�p�m�e�z�f=��	!�}���EY����W����� �˨p���	�)R�*��������9m�!� 0ݐ����M��X�J����+�X�w��O��?�����������󃪃���j�3���?c�)O��1��/������4h�-6���gM�fܼ�:�S��I-j]���v4�^;���/���[?�>�C��Kv�n(��MsFЃ[р9��tW�+�Yշ}ߏի_�K���]�fj���/k�����88���6=d@�)���yac�a ǞZ��M]��TJ鏽��g��)��X����y#J��Ş�0�]{H:��&~���,�8U}�Sw��<G9����I����!q�t:w�ܜ��@�;��@�V-�y���!����Sf�[��g,��6Ŏ8̤6k5�I�A��ib��?F�`�n�r���h@yc���(W>�3�Y��v�=̌4�;;��)��-Zf Ǫ�r�-g��� 8k>*2�ƓzY:���	�����ː%�<Gb�u����N�!���^��ut*����H`��2ᚻ�2cv�n��G��]!�)��I� f?(�J)C�X��8���@�3ݭQz��ib�:T���%�'�`���x�vm�mɪ�]3o^}�e�2����a�a����0����3">N�_+��C{��'G�ho�y��( �<KM�h#ާS��o�> S��9�'w`�c;"�sɣ$�Է)XH�}7t!�~����t��Cs��l.��&�n�z�����DxR��U&�@s�l��P(��k�~�`���
HS֞�56�����%e>}G������}x��Ox	��k~�m��?������B�r���[̆�g�.�|Kgl�,�ζ�3��N��2B�EC�gN�?��� h�:kE4a�6�jO�5����{l������
�{p3뗳�{��Q�TX�(�Q�$6P5Z�Sd88U�!0p����dS��v�;q��L��PP�!f�
l����Z��j9g��:�c�ج��|Pmq�Ӕ��g�|���m�Ҽ��ώh�y'А#��5X:"�Z���&^lכZ�׵\�a`�5_�%�������S�c���zU������{G��_���8~BU��'�L#���g먎̡�{SՆ)���4
U�N&�|R
�����߾Q�Ս���Z_�>�~ǧ~R]>^�R�]��ͧ�����=ur冷=�`]{�Ѻx�J-�.�V
��O��<����v!"��U3_�h;���)~ί��8&F��Л����x�&c��a�ɨI��<�+��eC#�w5ڜs����n��dHro����T���()�V7dz��e;��5�dR��g�����:;9��zMz�ŋ�Zp%�cK}	~�18}ۯިo���]?�3o�ۛY�/]����g� �Vf�"M�z�t��$����b)�`�0��nz��tS���pVkS��imO���/���>�Sꕿ�c�e���zAG(�p�}�]:'�yG!��K���j_�����}ӻ�{��O׿������B�/>�TdO�I�Ѕ�f��%����*N�s�k_VvTL0��~�^�9���L)(�mͣ��(-�A\eA:��kO�0��4ۑ<p��/�$#����nz�-��t�N#�;48�r�$C֑ө�P�t����'�Ѓ����;qN��K.���'�d�y����0y�{�O��ǚu���S)�у	MM:���!0mnk�%��;�c=����YO !9��l�PRCw�F�(�m\ӊ��G�L/W��^Ԙ�*�]r�ܽ^}q�ș���#���QLD�+�Xc}�Y^�ұ7J�~���dH�븏 C=�V�'���������l
2ؐ��}�MS�%䚰Ç���@�M�v>H��wL�N�ʓa6vv ?�J);CP�;���ZǾ{��# �G?���
P��Y��n]<�4G����,����9�4;#��\Wg�Ɲ����ѷ9�'z�m�	����KR���M�u�%� ��~8��	T�>����4�q��9��!Êk)m���Eĵަ ��\��1H���f5�r>#g;�` �	ҵYΜ2S�ϲ��6O,<�8�O�e��z�',?�[��?�����E��%��K�ϯ_�C��d����[dG�~L���ԛ�cS|,��tP��se���$΍=u�v�t�m�j*�h�5��S`�$�)����bX	����C}���̏�#�Oҩ����sę�p���);�;�%�T(�`�n�59��l3��Se�A�O��Ԑ�=C��tWdQ�� �{��U.�j>�n�f�hpIz�Ѐ}ID�6��s�4������n�DWo��X[��#�ZR��M=�R��%N)�/�����
�kW�\ݭ�\����s_Z���s�ɘެ���}w��/��n��t��=dN���m�C-@M\C.�gkC���s�]7�nC��D�!���I�mM�}w����'jw���ǎ��c_T����./j:������޺U�}׻��ݓz�����/zq^�(��SM���SB����ܱ�_;�I�W�1�.Jo~����Os 2\z���0�6�ݱ��dYd��1�J߻#�$^��Fd�==�4&���x����m���_�ACGJ�B��"u:Y۵�nNy�gi�kA�0D�@�)?���PC�P[|��m[t���:�x�γl���.���ͳ}�������W}c��M�Zu�@mj=]�lq�6���A%��YRg?��ˁ��t`e8˝X��ìL]߭��i-�w�?�������7�G��t���dHP����P*�\�ZFl*0O�vU�_�����_���7��������B�j^���Ϊ���q��"�k���r�mh:���$�UTa@�Skf��e�^�j��N�ѝJ�P�4�y�f�r��� �������Th�,u�M��94�9���v�r�*�Ј��}o!j:u�l&�ݠ,����D�'��ҍ���H@��iݛڧd
��C�k���8����CȮ�>�<#����nQg�΢������|�]��������ǆ(�g%Y:s<��g׵�U"_G�M[:1N� {	T�"ij<;3N�>�i�*fR��`U>�]i�d�t� 3�`i�F0�-�=�^&�j�Ϩ}����SY/����я68/ˡF�6-�<9{ȡ(���'�ZRӁ��d/r-ů�λP�h����zm����]7��n�A��rT�`��e�Q[o���\ʚ�}��#Gg2j�	��71<7q�Q���af�A���a��|�?�/4[� �ɘ�5kB�vCi$�]#��?�6�KƆ�� �������w��0rJYt�3�u�	p���M�fo��F+�yr@��$�؎?�x��ԑ�����01?O(���f��>�E��g����Mo�׽�u�A%�{y���J'��Z<{s�N����?�p��n���D�p^xjU)N8	�H���}ǜƨ�p�YN���ҽ�w�QIf���w�'�4���G(�9�E�����l��%�>
u���P��y ����%���鶖�YMד��u�����<m'jlt�����"���v�88``�*�+X�z��gHi�������}������ۺO�M�~�ˁ5���[rC'���4x��=��6�g`Om�j�]�b}�>�y��?�%�q�=w�iSdL�櫾����뻃:�aD���3�P��)�8��4~���@��bsVW�j�E�v�$(R(��Fpv����m��G/ԟ��JS=z�f�m�֫�u�V=�����?�����������sNO�R iCO�f�Y�A�iB±H<���e�f��@��v�M��ֹaR�\�\��6ڌ'R��Ð6�C�R��i�"D+A)Q� �ެ���Pu'�N��%�Fi�����C�x�X�s�dB�p�s	b�wt�=88`C*���t>�2��=�AIݜn>���i�x��:[�����t�
�)��#_l�@[��M��d}�7|s���U�����Yk��b��H��:�����#��%jW��{����D:��uu6ج{��U-봮���?������Q/�6!�D�E:�������c2�S�X��D�2� 3��uV��׾���;~����u6�X��q�j�z[���ƒA�ɉX��"#ޟA��H�׏v�Z��"ٱ�V��Cc`m��28�}��3����c�U�bf�Ʃb�,��<'S֛�tg:S}�QnT�����b� z	���(q9t
��аB ^g�`�:7�7���F&=ߞf������g�G'6� �ns 6��S%0�.�f۳�퐌W��S%�;k2��s��8�C�g[����/�mC�ЃJ��OgJ���s�C�)��m���}�g
uҺ��%3��{������Y/��dS���a2iځh����}sMl=�mp���  �k�nDH�Ҏ����	gqVs��B���Oݴ��A>{?�z��w���}�����~Cs�L(RVW����~(���f24j�@��y��z ���Գ�!NT���3hn�u�L�E�҂!�L�H=�+���@�=��D�A�?�>�����e���6�6�A[�C����B�4������:IQ��Ɏ,�`:��~����{���H�VS�PZ����������e��u&��7��al�J��6*�����%\���5�
?l�>��������������t��3AiRӋ���.1�FS��	��<3)	t����@�������	�m�D�\dx�s����oڳ������pd>��9�g�1�Au7�h`��G�aK��n��,�l'���?6���9=�ѣ��c�;E��(9��]yg����|7��nV�����Q�����Ϛ�wvRg��5��U�N�)�9@I��`��N����'�4�k����5J����t7}���L$l�ϡ`O�	j��>-�7r�c����}�e��ݠo��'�=ӳ����G<0���>�C֘>G���O�F��U�Y?��ԍ�6P��m�ͥ�z Q� �Θ2:N�
��{Jٵ*�L<�K�y��
�)޻Q��������_����O�<v��/�Q=�}��5�-��Cׅ�W�ݱ�"g��U4�w25�G����)5(G<���6k�s�ʄ.r�;O����K!uD�u(�����섎ڸ�X$�S��C��hV7�������i	S��10��%i��� jD�������é���@O�'K� "@ݿ����t��J�7P`n0���C��� L�Z,jyxP�G��m��    IDAT�ਖ�G5_��Y�r3�A�eA��}�zݾu���\��<P��a�y���KfY��UսM���7����o�_}������s�f��y:8;( 2��Ί#�%*%�� ���ۜ�~s��:��~�+�K~�gփG�f�$o�@�>��w(��N�c��Э�x��O���5ozWݛ^���"��!��TC̿��޾2�/�i6�Nj��h29	F�U�f��3-0��,~dK@��%N�p�ֈ�b� �i!}�*;'��;n��)B��k�q\�9i�"�rʈ8�s�b����f��K�s>s���9H��7r��Q7�q�_�����5mq.9�~�8�I�)
j��,�yUFNH+�!7���7�c��l9���]�q�[�B��u@6��Q�g��ͱ9-����~nN��%�l��x�������G��������������ʈ��3����d�L���9�Jͽ�,��\���'~��Z�
dZԹ��d-�|��䚚��c<�K����H�3P%*w�Kr��l~�@�T�8�^}eF+�΍$O���g�@�r�SpVt2�z�j,�m� ��F����9���[���d�ީZ�K`قw�匜[GSD��;��䰿"���k�5�v��#�2�����GYRP����7��
�C�vcם�	��ø��i����Po� k�N���x�ډ��!�&8�`` ����0����V.��f 4=`:j�BA����_r�F�
d�v����O���L�������o|k�7 ��\�ˬA�G���ڎ}<:;@�N�m u։泳�z�P���A��(������Zr%���x�l����y밖W��&I���1�;ݧ�e�:����J��~0؀���s8������@�$�!{�ϛ	
�l���G�l��)~��Q����1n�%��ֻm�n��d���rZ�Y18ő�ə-�?ʷ�������-�S��6�g�`،���tb`dE�y����|3���Jv^`o�K�����r��H+1�}�1l���l���K4?Z��~�W�:��fh~�7��;�߿�ucs�#4��m*��{S4mG��5��V��H�K2b|A2��� �x�_��t{Z��O���������U�K��k�u����rZ�{��'��ӳu=���˦�R*�`0�;
t�պv�um���@W���n�_sLʌ*S�C�#A��
Ep�i����5�ɚ��$k�\o(���ʚ<Jo-'&���2�LӔ���K���Wo]%���4tP���'WG2g(ǚ0�v#L%���i��{����g����z��nK��h�gP��  d��<��.��K�����(�|M)8<�³��u��:9�S/_������tSz�`݀���T}�w�������z���lzX����7E�;Y�0�u��D4�}L����"(�?�W'켻��kz��<�����Z_�y�Q�\�A��B�`�������e�~��g=�jc�Qp�z��z��o��~շ��y���.���rmRM�5[�j�:@��8��]{�0|�>�(,rMj�M��F3SjS4_d����,ސy��6��kn��c�L�5��?A#�F�򂐮��c?`�7���) �s.���]���{F#g���MjiyU�Y;��.c��w��W� ��f
=�8:�����}<��Mph�S� ��x�.��3��W|f�4�`��s��6$�$�:6k2�ǷlH6-Ɏ�.vL�r�x=��Ձ#6wZߥ9���ʸ�1��.َ�l2�D��#s`mt�@�z���P�#j��W�X�:��_�7�d�1i�A`W��
~��=�>;|rj�18�9�����9l��C�j| ݬ%���q�LgL �qzms��J㳪��Q��{.��� o�C-%1Nϙ��N���o>K7���%�ڬ�wCO&�Hc�mT��7�/5 B��Yת�e@���h~w_�1��>n��#�萻��t��A�pϷ�I�ϒo��5��ut�v�S�[�`<�`[d7��7�����{e��,�f���7��β���ғ9@�c. ��J�����}�l�_��"�##��mH��^�d�(3�����<zĲ���	��1q
 ĸ����z�ڕ���z%��׽�������)�D7�������8 �?�B�-��ՁԀ,�3-���NuQ��O�5�J�~O��YYkhZƼ���<P� }��t����;P��
	ؐ�����~"�#��P�o�X=aCM�|*y5���g�'8��	Ҿf��y_��6k��LP�;�􂒦��[���V�M�jàt��0o��fb�b���8�>��թj +®��
>{������9�6�D7'l�]&�6d.FG�ǓhL9�Az�R�3��4^��֧�\ߩ�������>��ʘn�����ӿ���~�-O(c
%�����t��,��j��T2�NYH�+�MX��ô���y���|^�ӳ�U=�]G�{�Q/z�>�/�/��W��^��Nj6����n�~���w�x�Ѻp�5i�&	��t�����:�w��P���ﾘ3��F:�R_�nh�|TQC=�{�hg��_���J�B,qΈ Ek��������k��^�C"Z���l��s-�PqkRIA��Oge��fLr0����ɉ#؛���J�>���~}'22)ؗc>:2ڢ+��A˩8���Q@W�VW�Z�dQ!��!kz�έ:>>�KW�T�t�o+�}��V?u�����������n�k3�\GW��l��SU���Ԗ����\� D�5�lv����b]��	3���{��|�g�~��#W� �)IIc�c�^�n#3�ez�#�0�U��&�a��8�W�̛>P�}{��O������zV��kΉ��ȡ[��8��l(1�H�-�u%|���4��-⹴v�,(á��P��l癊C�u�����T��	'����<@�����D*M�����r�ݱn��4nUdL[��p���ub򙇔����$����a�0�JROAW�3����5�>���@��E殷���ܡ�q���-=� �g�N/�3���4B��	�耄)oMǸ<�����T��;�4:�	���J6u�Qg�$HI�RQx�5&��<k���7�S�Œ�����w)��=$hߥ�Eu�t�htT@i�7 �@�L 4�Т��V�|��&��c���?y�0�`{W�{��������,b5ʠ��t9�7�'�mo�P��r�t��Nh6�"y�q,�k�)���	���9Jn?�'l��5�~��le�owRo��OU_&��;u�EU�J�m�[�������߁�f�/F�;@�� ����L�\�d� a��ą��ZDSI�K�5\�@��-������>�	k>SL��oh5���e�t����5qC�W�v��r�g�&8K�z���%K�3�iGx������o�f���]r?�h6��#_�O�-�����oW��Mo��՚ <�vQݻ��O�>����j���H��HS���0�b��FG�f*IHY�8�_�z�Aa^+߬�q~�h.� �C�W��z�6�k���1n����zZ(S*�г�/q��`f(�Ldy����l3�(}S`C�.����VsŬ)��,C�	�׳mM���#H��f�u<s(�+��A� ��8�*�PS�!��L���D�}2��=w���k�r��t����8@5��495�nFc2t9¬N�ih���9O���i-�n�K\�?���^���kL�C`�׿�;���D���
a%�$��[��rmnJ����Ѫ-��Hܜ5���c=b������w��-��G.��K���?���Ӛ��xwV�=�{�oԍ'��������j��=(|�+�\�=ҳ�:�}������q���3 cC��M���\$�{D�U�?��l�� 4�Dy�P:�݌�3T2�C���,j��xپ:%GD���o�67c�n.zQ�4Z� �a�^��c��ϖ��F@7,ɠ p�FA�H�Y�c�: f��ɗh��Rs,8RJ�\Jd��Ǻ��u���z��G���E&"�ӣ�f]7�?Y��I]�tQv���{�2�o�cd&�����C?����?��z���^����Ύ�Pf���#����FkgJh�\A�eE���d����''��ݮ?���Q_�E�Y����b/y:������<W`�ܦt�����xA����^3v�Ep��^�����������^������Y-��;v,Uv���F���(Qd��*���^�w�������o M�3m�M�3�@YQ�x%����]ch�4/wO=��"�OnP�4��쑱�ƀ[ĵ�tP�,N���9�E�:�3�=՜�0S��g��5�1�����^v�CF#
E��l�Uۣ��K+x�K�2�t�쇉) ]�9uJ��.�r]�Ԇ�F��s:�� ��k5�vB��}� �N�T<Z��&.Z�w�?L�Z�i�!�#$�Uz.Hu�us�5 �`C���NZt���V�$0U����H���:��e��Ph6��Le>;葰r�P�dOT��;�&u��Fԍ��YS'=0M����m�g��a��EOz����K��Ӕ��ґ$j\įvS90��h�;o����)%�S>֟I.$� ���d&0��I��SR^��ڎ��r{��Иi�[�.�[�.��"q"ߠ:�Ӳ�;����H�94̮���J��6�<����K��@�1�+&�@�e�|��q���>u/��"�rv�38Pe�d���X<Z �`�Qr_�\Z'���G%�R�rf���͸�zd4�dW����#Ջ_�|RyoܺS?��Pg���;�D>Q�V�2D�¶Bs����Ȁj Y� �d�'���Z9[��b��lc,'9�_R{�E���a�� ���#�~�����>��|��>YϬ;Ɩ��R� C�����!����1��b�~(��yR�}�gԊ�� Ug�"`+]�����2#����lj��l��}MS�-M[�#d4�����mVgd!!��C)�sL3��n�&PG55ʹu�˲�ףcƹ~�8��#�8����kק5?�U/{���W}Y�쑃v��y"=I����|z_�׾���5o{���Q��q]Q�Pԩs�F(e'F)�n��X�S��Z٫����9�@��Nk�����f}��u��?�G�N{�]3!ZnW���>^�ժ�\{�.=��)��w�n��۷nԝ�7j�Cpt�w3�\p!������#<Lb��)T����um)��W�ʢ�����Ҡ���!M���BSv��t��7���p���9-
6�q�Z�'�	8�eß�is.s�5e�IgC�N�o2"`C�9�,i5A���.��V��r�/׵���+Wk�<�B�9�Ҷ����{�	f,/=p��:ۖ*�$%È ��{�^�so��G`vwV�%��Z���#�)k+TP��4&3�*N5ۚ�����:^��xv�>�?�����z�K~^�R��h�E�ϗM�=�����k�<֕p�:���B��N'��ݪW}�Է��/Խ�ժ�����5�y�����g�����n���ON�P!��0��صԴ2���߬V�!��ڝ��j6�i�����<90��t���?�8 �v���5���7P%��Nz�]�`�Q�>���A����qzS�`�0��F;΢W5n4��;���
]�� �v�7o���)�M��H�/�F�w5�1]����;����!b��dE�ΥF:��ٓ�e| 	RȮ�LW4����p-p#��N��,R(g�IӂC�%Ͳ�ӥ�/e��	���L)�R3f�7g��dm2'̘8��dp ��v+pS4Q����C�l��p_���m��2���ſ���6����^T��n�wE�Q���Ԅ��=�MP���@��wFh���ॴ� �=�KE�j���FݩμS{��t���������HF�ug���t� y��~e��wH�?�v 6�9�H=�r�n��閆I��Qw�K�Z=d=��}'`�{7v�U�8s�$�F��� �샠�@v4�B��@oG
7�V�jk6Ԝ#Q�:��n�� �_� �k:����z��̌���NBAI阁=P��}��b�ޣ��-m`�ɜ!��1��,\�	 �I�n�lL�:�P�Y>�_�A��2����G��-[�|bZ�}�ם��Z���(���7��f�L'�X�fP�$,�/��:8������9�����f�<c�'��A>Hڃ��/�T��B3�����n[�ɤV/2����¶��D�Κ{�p<�}�'���Ld�����Z#��w'-��?q���gqs�"�$� ��1mz(�@Ĕj��7~�duR�ӛ���;����/��zhYGC�Q�O�����&L�������_y��M��u~X>\+��'A����-#xx�H�\PHI�Ŧ�s���'3U��[�ñqV�59�[���W�������W�j�
bh�u�n]��ן���x���ő靚��;7���u��m���+��;�i�b����E�ᆳ!��Jh ����hЁf��������3�@�N��d�Hɛ����lѩsCA��!$u�|�3�#=[��7������C�chǹԛ�#�����dR�qTk��Xlݛt��y�X�05Y�RtnT?YF���p*3МJGI�=�<6Ò!����~��޺ɚ���W�����R;�������t�_�;��^������B��&մbȤ�)W`ʚ�A�� ̻�ƃ��gu4�[/�ן�#_X�Ᏺ�.�Jb=���)��sY�ޏ1����~vp�d����5~;v"������?}m��ƬV��u�_2kL��4�C��3E
JU� e�Z�縐��Q]L�s7\g]ym(���I �}�M"b8�<���2!Q�tHM2t6X�CJ��I&i"��s�;�}FTQQ9�Ԫ#�2p�|�2�����-YS����'ʈZ�U�]bq������^|�q�P(9��5�����M_�B��	j1���z�)7&@�w��J6wH�i@�����n�Wk
�JsHc< ����z�?��@f#(Gr��Xj'=���_	T�x����}]�ˠ����>N���;��]Xր=�#���h	;0 �=�g�|'V�C�ڱ�Du��p
�LN��-%[���:J���()<���� �k�W0�u�m�v и�T�Ն,Q�7�\�-E����V�UJt�7G��c��C?��T)�*�� 4���ɁjQ�M��6Ю�F7�Q�٧ ����>3К
���}��qǳy��4�s;@h�d��y����,�דe>cV9� �<-RTv+s���~�>~'�x?�1� H`y�6%�}.ݜw(�-��Tn�n��|��`6C�=�1�msSP٫PAm��Vԯ�a�@~6m�40��B�~��J�뀁��%�����>�-;/T�M��f_�1�Z��kp>y V�u]d�mn�>m��<���I�v��� 1��M�֬՞[K.�1KI�=�G 0��I٬H�W'���@�~	)�́�WȌ�91t<�|}*/�p��X2d/(!��,�D�����!�/N�XMvuo�a��n_g�m��0�F��ܲWl�iĎ	�Ae1f@�f`�J՘�ɩgqH>%é����^z�es���8B)�����HĬ<������f}��/����/��^[���;
H˘>����_�-�ӿ�dݛ]T})��s�����urTt�����9]HE�A*�:&��ș������Q��٭�k}��:�ݪ?�ǿ���K~o]@�]�n�rgw�΍'��䤎/?X�W�U�(f96uz�Nݾ�t�ݻ#E��2�s�|��~���DY�Mz/�-	:�#��4��A�]�3T��>: �GWg5�$� �\	�ZAGy����f�9�g ������\�3X8�EYhV4 v���c��u�s�:�����l��v�A����]�G�9R(2^��I�<��Եͭ�k�4u����/^��{A͗�rb�T�����'�����p    IDATu�ڃutQw�8(�P��'��c���7���W����7�fǏ���J��B,@�����)D��JB�=3�{7�����n=x��?��_\��鯨92� p���٨�@�i�6׳��4�s���/����� +�Bn��{~�]�w^�mus}�5�;�3i"��L�����O�{:�`���&�D�U��j<v]E���Y�{�`�"�����s�� �1r+u��D8�x��:�|t@����t�K8�h3[��#�`��1�x�\IKbf@�\�~8K��|.N�x��Iɸe��1�,��nt�]�@��S���^����ڠ��r?��J�{:b`�[�%��� ��qJW�8�;|"��4)F�]R�@��f�� �Y35�J���9����5F�٬)g���8 g���`�Rw![�㟚�o�_�8Y28ܬQ�b�ZU�6>2�vTsJ$܎�a��.AёH���cJ&�ЍN�K�r�z� H��g���I`�h�!�V�:TR^ý%�'�#g��J 
AR+��u�|�А=_��C:8'{���M��P�)k�1tɌ���f.�D��}%�Jp�iemCIiC@�޺���9����\���I�f���2��j3�w�od�w̝d,���\?l�:���^�>ѥ
P��Y/�z�!Ћ����KB3f�9Ǝ���<�������ݍ7ǽ~>��=�n�CL}��t��� ��u��۷!(�Ttr���FJ.�h}�̢b��j7	��GI�f[��Oꉛ�Iv�L��1'p#(��g�`�Y�˛�Q��mZo�����yJ�ΔL��Nрfg����}�7сX�5�YHJOR){f^�(��ԓ��D����UBΞ�gRTt���,@_��;��5'�(1]��"aJ�7FpEc�Vtم!������im&�Z���g��Z3@u��nR�5��짡`=`sZYc�-;����������#��׭���sFs��_�<f�Ȧ�G�4J`�����>�[����]����1]��1u�5��� 0����wި�u��R�zX$� ]S��SQ�Z��bV��9��x��۵A�4�u-'ۺt4�����oO�pI����`~XK�yD̽�w�u�w��.O����X���������IZ���[u����/\~��U'�H����³�t_��z�� �Kt�nu�c�Bl �1�Xh�9;ֻ�W
�U��\H�k6L���#f�4:ѥ��n�	�Z�
Ĉ؛���?;�B�#gR:z��TzW��eVW���
�u�~\�"��� Dn�A��dg�[��J�]��VFg@��q�oB��n�E�����l�I��<ˆ��Y]�\W�=̣f5M�uv�f=�ws]/_y��ˣ����c��Y��O+V����?^_���v�v~�&�cw�5���D�F���3�0� �f[�[�ٿ���+����_;d����|Iy�[{��??0YhmC[-/�h��ޛU�뿻��O�����T@�)�@���s���
�:I��Be7${��]�-$я��<P�~Q�Ԅ
J����F��z�tT�3���%���M)�LK�����ܨL�ݛ�Ր�{Ċ��Y[o��m�Η�4��Drmw��0�pf!� ��ouRX�nlv��M��qI8-C�jݵ3�c��<k֔��"�SS�Y���P�.�	���ԡ�)��^�0s�ls8u�׿�����
��w�p�]��:�-@bh�A�3�(To�^�6&�k���X� �H���������cB��*k�h�,�p�Li�~ks���^pm�k���.������e�����
ȘI�o�2\�CӍ ���Z�k;��e+�e�hs-�pyg��=v���8�g����zlt�e�R�m�4�-LGm
l�&��[��������gZ$�X�/F�s<�w ;��K˙�'��c+V��a-fn:��|�d�(hNF�Ԙ��s+�I��۽��������7����1!�e�D]3�q;-���4�
�~N����iN�XI��� #fx�
��K,A&vu�w! ��bA��[����~�����!>DG*{��&Z��&5dS�s~�3��M�?W�� `��<;;�9��I�m��k����(��F<�P���Ӏ��T����{�86Ή�5����0�jW�_Dw{+?��T'� �d�e���&VȘn��g+�e� }��h�3��ėh���M�N���\����]�MM�	1Li�ܽ���{�ho!�������q�������(9����h[�%�1H���ܚE�� ���53�ӓ���^����m}�ʘ�S��՘���������䨶�ym0!.�j���6g5]ݭ_=�O��Wԇ����8�T����������Ok��W/y�������z��a��ܩw������}C���{5�_�=�i��~�ַ���'�Y���?�ڿZ/}�c�߭Ĳ\�ֽ[���.t><��ϖda��nݼ^�wo�|Ӊ��r�18�B"�^�k���8�BoT[
Gtyp�l�fI�&O7�����
b�9n]���^$XO,�Z�4��@H(;�B &�9������GR�q�b�f :*�9y��]0Y�#����\�����<ͧ�1�����t�4�h��B�s4��q�B�q���ge�&u|�2둗G�*bߞ�{��y��W�����!(�Z�=LG��j��֛��D�������a��krx�U5w��.$�pә��)���1�% "zZ�:���S�����W��z�'}D�����6*ɖ�Nc������`i�����z�����G�\��@��_����˦�M�Yed(�;�v6�D�L��Sb�jt�GPٸr*L;'��;�*8�Q�3@&RwG�'`3��:�kK�$00��fP�}�C��.f˖9��g��:$�����m��n�����,��Լp_���5���Yd��}1I����'{!T;���)�=� ��|j�Mәl���4%�u�NwZּJfd+;�`C�8QF�U�������C�f�ÑW�a�c�<�	b�����p%z�<�Z��NB)]�FE��֑�gԑ̵i�lALzcn�P�|~����^�}�сprҷa�	����f;k�Y�����ҍ����F_7-�=_G�-�ө�
TJc��;�`F�ig��~R�Á3��=æ�#w�:L����sx��@�hs�O۽n[;��ex󰦫*ؖ>�Q<���@ Xe��8�OV���XtF9�a�&qȭ|L�MB�p�z4���ެa^�II;�g��~HS�֙-�h�d�e���C�)ku��N�I�T�ٰ S��:�.���<s��1� �;4�n���������bc�4�,d�a��9�J��2�kĜ�8�F9�[��&2�y�(���!\�m]�r�����;urrZK$�4�
#���O|Ug�;0��ӯc��]x�w��/��38�;I��濹_  g|~�Z�����ɭ1��.h� �\�?����~1i�P�ѹ;��Tn��dZ���.�HO�Vp~n��Jj�TӋK!�T3@R�@ߝ��k����p���-��im.>_kWk̛�3쫓�S�w�%�,��ҵGjy�Z�'�Z�f.&}VT��vù�وL�Z{�n�d�T,9�����B��[Gt5�%�K�y�n��K��������zŋ�00}�K��������w��~���dz\k����/8�h���vu���V��_�;��~�'���;�U_�O�~�G��5����z�K_X�����/D�Wu�n���O����k꽏߮�z��]���Suv��5��x}��}Z����g�klx��G�\��ٚ�g.�>���Vqȭ[7Z2����cdB�⹙keIHg�a����Nh�M����ڰ����P��������Bu��RJ�y�R�+s��$�_݂e4Հ
�L|>5���F9��e�@�%z��FI�"�fH����d�T�"�lt��Si��T�%��h�gO�k:U �A��j�N�9�t"�\�����dRG/֕k���������?�D]�x���P-/^��l�F_{���i���U������W����.���*�u@˴��;;o�J�&��ʻ��OOjr�D��^R�/����������]��s�3 T<����9�� ��@	F}�Z��w�w���׼�u2�Pk���@1���t7S��7&���\,G�s #H��D�����9�����{��Gf�<��*
�mˡ� ��s�o{Z�����]�9S�t����X�
J4�B�	Ŏ�J�_bK�D��@Tzc�c�h�N��^��3� SΔs�9��~�S�����������N�{���_y��>����eB�wf4��*o&�D�ٟXQYVKU������`(�4��N����f�ш{~>�@�Ԩ�P���O�%�1���6��ӣ��}�4�T�-�b��Ӛz���S�5M��VLa���?wr�+b�f��V���v��@��\� ��#��
�,�TMm��9�H��W�� �@Ɂ��(�O���R��$$����L�r!'U���`�v9f���Q,��Q$hK�SPd��zFKO:�/I
��b.���>�9��	��bږ��J�Z�Rb-�V�D�2g�����~/��Ά���b����Ɏi�*��@���*�2(����ML����]Q-��߻P�<���( O0B�_�| ��`�U�JL}�*(^y�y�5���4@3�AI���b<��Ý?Yp�O����J�׾� 0��mSt%�$��P,q_~�����7Q�Z[s�a�&�&�qv;���y�xx�BG��ͪ�_�KF�q';����Y�^�w�'��;�v�+�By�O����T�X�*�h�/(����;>M��E,��R����~p\�����{O�������|�%O��Y�n|��<��P &�7���V�\2V<�R�.bΆ	aA;�1��[U������V�nd���dT�K�D�j�nCi�uk�D_��R�pȶH x��:�;D�l>P���@�aŔS����NakD?�� .�����ye�g9���&�� �P?�l!����hgg'v��c�h�ŷ�ƹ���4�1�g�@s��QI8c�b�LHQ�ʼ [�ض�d۷��ב�L��w�W��-��z U�y �j�����3f{�r:����������yA<��~F��91�*oVL���u6�c���^'�L�:�It�{񅏼2~�۟�7Ac�����_����¯��'Oc�˵W^�}Ɨ�{I�G���9�_}���w�����A��˘l���>�M�/}A<�9O��0��r3��u2v�b��޾A�77�?�������3�š�����Ӄ�B�A@@���J��ɩi���Y-�_0@R�J��2K��鸡2�N���"<��Ƒ�YW'�X���B߭M�8��攣GԽ>����K5NԬ�
��T^>[: '���J�̰"��j�`Ȼ����Q��w�g�0�}P�V�+�J�a�b�Rw#Gϟ�J�t@R����vb����I4�ԩ{���'�7����ZRtS,��i&���,;������'���b�Fw0D0��n*C'�Tk�f:�<w�e���Yn������yQ|����;��[e������h��e~�/F����r߉<Ri?"��;7�/��ǉ�ALb�L�1�U#\����K5^��PK�	k8�c�@`[�I���9�:3X�3D;pq�?���7H���,��P-%%�NtS�}m��I�?������iF����Π��zQ�Ʀ�B@I쫪���C0@�h�W�^7�#&WQp���+�ʯ��K��љG]�!湭D�ICF�8�7�w�Ι��N:��!��=x��;�Ε,�xE����QJ[d@��v�Νz�]1E���C�D=�x�G�h��I���L	�y�-W۸�����P�ݿ�Y����]wR�"�U+%�|V����A�Q��s�J��A���O^uVs)ڦ�V}�JF}ku��-�`Ϟv� P>�L���ǜ	-_�>eX�&�>��*�Ĩq��"	T';�O��5p}8W`P��ő�r]��A1ɼ	x��8{�q[P��Z*�j��e K!� *KIƻSm��{��B谟����c�"�i���Z0%GM0ր�OVOVxȣF嶝�sk�
��$?��Np^lEs.`SZ;BA�
���r��?�9ʢj<VM�[�n���"i��L����(UQ�uM"m�AȜl5c%2T�I�4�j�~3�s��Ib�_{u<�kbwo7��θ�O�2������s�dO![O��I4*�.���<�����|�����_ҿ��)�«rJ�9Z6b��0UP¶�S�������Ŕ�G��g�H\6�Y�7�`��AjF�����LG�a.�(ע�B�HE��&+�� )��C�Iv7���X�4��;]�	Ві���Ǚ���D�)�d��c{{;���8sf�h�����mF60SP�Oٶ1�i.0���.�tb1$������"JJXi�1 S��� 9�m�e&�H����Kv��t��ߋ]�/�?�k*�h�������������__1ubz_&�7��x��[��]Gb��<J���\��rGz���g=%��e��.+*)�~��;�����;��Yƹ���'=:����a\z|�uz����x���x�{n���$��'�?݊G\yN|��__������ a��M���������egO`��޾��V��!������ Q��O
B&d��5}V@�ч�V804]3>��b��$s:��rc$G��Υ�u81���\��$UYtУ�)*���ұӉ�,YUU!�-��ؘʰ��G�=��|�tHLL�LRn�E��(�,��ws�$�S��+Zm�>��⹰�D��z:�2��0.9J[�.�:!�@3�J@c���S{{����� Fk�8~�E��y4���XAy3��9j�t��|���џ����m[��8�^һ�XC�)�.�8p�s-�*u�g�]�F����+⇾�EqŅ�T�&&�h�:Z#��ş�������Ɗ��=g���, E�z~_�����e������y̺G�h�whN�!�tf�&��$	������:$5T�)�>�n:l��VT&�H�������;���|��"�)�clC*�G1X�`m�ѐ�����yG�p����U��3�@��M`�3�$�U2T��
��O)�P�g��+'jp��r7��XO��k�0� �>�o,e�K�+�(�D�rX���rUB�G���f��'��P��u-l�C̓��ժ]��#y�����t%FeQ8�~�,4��)<���V���$����5Y5=����5�E\���SNnYi�]�}Pr���qE����3�$�����f6�!L���^��Cpj���TsOr���fe`��� .���~7�AI,x�>��#ft)�Z���8�iV'�&�|Y�������g�}<$X{�=�����e�+N���w�b]�~Uj�yC�$�J@���	�!�Ӡ'��l�2�-�o
5:�f��:L�PA�$ʤ�Mtz#�hF]���
Z	ЖM�7�ӕ�
jWК'�TL�d2isB��i�Z~|{
iL�- 6�X�"N9�ǔ��19����2cRT�q��Y+��ʟ&�ϭ�U�p����N�~9�r9�Ĩ���~P\w̓a��;����qfo�^&�d�~�Z����\
�51-�y�n�E���|i\��,��_��;�u6 H�Ap�` �;G�-��]C�n[�Y��;eSl|�����=�@��	�ȘQ�$;�v�6��c�~���w+�\�n��31�;e	�7ch�$�/�W�>T��W�)�v1��,���
0N3�[A�7�L%踳�'�'Μ>�`+�k��Gw���f�l���2k�����겦C�HC����wMA��QXsU�(����|�bͳć�F��g])ghSym�3��3Ovc}yOx����oxj\u���Tu��h�i��� $@ۿ#~��_Fb���F7�w�y ��$�9>�����    IDAT���9(�f5�7~��s��{b���]N�ӛ��~�C�;��������F,#n�7�߼�M�'��8�ލ����ً/{������x��WD,'0������jh��H��~��t�F"&Zi����0s��d�>S;��)sd��N����bt�ih��)?C��{�%���B�En>�6����*m�cr�)�-�:N�L�����:������3��֨e����L�iT�lX�6蘓ƚTgQPT Y���˒�*�GA;��foߐ��\iU�5�Ec������0Ar�#��V<���d/N�| �l��T����Kbcs3�kk��#:���O�*f�~�8������{o� �Y'�ƌc8�b3�CE, w�cG�'����L���ċ��U����8��
��ڷc���${o��C��o�?_	�4��	N���\w: �N�#�ٿ��������9���ET�����A*=��d1�E�&��jF�@���:��$�Y�%	��?�I�ERD:�J���4�dK��B":�܈��8��L�S� QI~}�3��?�`�h!���< HQTVD!�*a�5ׇc8�ۺ;�a �H5`���+'D���O5a��Ĵ(Ţ­�8t�Ş�%=���vN%$��p�_�4�����l�m��D���0}N'ժ��cX�G�+���%�W�`�v	�C(G�c���m�ϳk�@ ��UA�ڃ�D��n��\�P��@�[*}��5�g0��G\��^(ݩv�}��2
�G�~5>�G����BeF�1�z��O%���E<�
�XkPC���!Q{��3Oӌc�Mb>�� $��b4UJ�����{�5c N�
yj�*h��ha
"T��ET��{Ȼ��+:�����`e�T⪯�~J�%s ����A��T��X"g��t $3��;�R%�~�F�V"ǧ�-�vp�����D�W�4�$W<��3�ʯ+U����j`����떺��.�T|���0��i�k���.��B��>Mޛ�+��>Av�#�`�Ӄ)���� ��e<��+�sq-(���<������3��ƲfGi�u����u��v�w�����U��5��yn�{:9�=�d�z�޹�������o���l?֎���!�\�x(9l�I�{�^o@�G��m�O����XT�V�YL��~ݛy�{�ʫcR��Y�"�7a�!r�nz��iU�՗=�d�tWR3��}�u?&���:y:�lm�dol�U����?ڌ�ڑ�FT����d���*_����Φ�U,瓉4r�@j "3l8ǖ��ؒ���j�}�A#Hg�~U	<�0_�`'֗����<~�E_W�d�_��z�i������ig-&��H�ρߓ�xܵ�?}���g_��7܍��~�o�k_��8��~������%�������g=%����_t⎭���5���������'�������x������.�Q;;[h4�3a	�*����@ѶK<��S���� �P�ͤT<�N'F�1)�"╿;��d�UV�\j�Jn:�nI�&go*��p(�����t�m'��-�����%���*�{A�d<R�d�͊��*��5��d�Ri*b��Jψ��'�sEY�LJ�0�� �έ9�)8.S��q��O� QAQ�^FE*�<y2N�:t��/�#ǎ���z����e�9�ղ��(v�?�������0f�c��oD��b���YeC�^�X���_"e��<ۊK���?}���	�yHaa�LM�*W���T���Kb����531�]E��M���~w�.�Ū3�y�T4n{�4��=�*�y��s)z��aJU?:�A��/k��%f@�s�^,3!͊_�Y*~'�*i,���b��f�ǃ��B14���%�?�(o�(8V7��Tu�R��T�+�+��=����&�N썶��)��t��`�I�_KI��C��~L�H�Jq��ʖ��G���	,S��k����z<�N�N���<��� �(��;���T��jʤ;n��g)%&[��]%��+�"�`����#e��}1�^7��xAg�IM��zS�ʅg4՛�~r'�U�(}��.%l�{*j�|��7�_���)O�Φ�x.�WfD�
u�2aeE�n���Sz>��%	 ������>T��הSgڡϝ+L���ojκ�8/5Q�W<���{��۲R�*D�t�G�E̪���LH������G��&�>+�q'_�eϑ�IR�^P�ªZb�u�E�)g�����bm�'8�c���L*p%��:�Y����rV�o��>g���S���]�	��gݭzn_kⱒ��^_�*hKUl5�|�
�Q@(.0�m���P� |-}�
 X��t��t��2���x<�Wk�\/����ĩ3�\�z��z�jb
0 �ұ��X'�*����ʓ��|��񳔓[@����,G�W���
I�'簞m���q�'�F��q���i��I��9�z�>�I r���b���s��H(=̵���Ș 6ɬ��_ A�k��ą��Ƹ<��b�iVT�)��,��U�|����$&{{1�݉��������vsv�Z�F9Ab�>|���5����	h��� ��99�sN�hN$k��g\\�4E8���	g�ɴ�_;
�c:i��=���X[��=���~u\}Lk�"�N����+�s���S�k1ˍ���j��4�vc�܍/�����ozV<�5,p�?����ߊ�ӳX흉�t�9.������x�Ӟ�>��*�֓?�c?�����,�[w����{����_��X�Y8���ӧc=����،t���#��cT�")�L���|"U,T����U;�xAs��?(w����Ǿ��@�rY)�	�����n�W$F;Hy/��D���C���B�u�4��.����u¹!�ˤ_ې�	"��x,|���*�bH��\9786�3�Ʌ���*H��}��;K���UՓV�FۤUS�T�z:�\^�.��I�|������3gr��F�s�9q�ؑ�Sm6����u���9S��;o��z��`u$���֣�3�X�6(h�#��j��A��g�Q��W|���JD�$W�iM��8�P�MJ�Jg'��>ӟ򻓛�̈7��M��_���[��e?R�!��`�P�%�AW5�pIe��\L��"��R��f���7"Y@�|��͂�:;b5��d�X�RZ`������c�����*i��Mq��vw��ɒ X��؞Ci�BVU�3mP�K�J)�@S�i~��3-�����D��wbZ�wNNL�B[+ �\��[����D ��i1����Ʃ��}�S�ⰤXX������ȢixN��:�ni�N��j�
���=�%�A�#��f�</5eHr��3��S��\����Wְ\Z:g�z���tU%�m��g�E�u8�	Μ�ǠūRQy���T�Ė��Y�g�g��*_�`�f����)ӷ��1�e|ݚ�;�K����n`���?�ͳL+U��Ew~E���1�<������("�ׯe��՜���
g�2PvEX{nZ�b
� �J`�
�dz1�v�]���61���1�l���6��v+�CdG0�q�A��J|nմ8D�n�e�!< WT�FO���?�I36��a��&Ȥn�~�E��fM��2* M����J?(���X�1�~��ѻ7	/^���J/��<�L��(ōI�_7�1t���΍��5����~GLgi��k,�d�y�F����΃e�x��h9D�����&��[M�V������BQ%�>�#j՟��~h��Ef��w�\�f$�m����-@��t������m�,F��R[L~�>�h��+1��"�i��̷r�J�W�����*H���X���ڌ�H:����ӱ�ߍ��$��<���GCb�c5bj
�-�nO���.�<��%�#�#�cOE��#m�?�iXq)�;��ĵ@�@�G`���s*�>!)7��UK��fb��G\?�⯍��P��3�����E���񮏝��n*oz�w�,��to/��f��k���^�u�Y��#�N�?��ƫ^�����O�����,bcs��Q��7��9�G?�ho��O��~����w�7V{�'��+Ϗx���}��b�����8�ߏ�3ۚ=�`Ӵ��"x(:0~�Vp\%@�1ď21�T�����م���g�?�7���Ue�0��NLyl�*���X��L�A���HRg��Ic��'��(|��Rii�Pp��՞18�ߧap�F�_ �����z�,�]*L���[�R������iLesl�Y-Mj���3��E_�49�V@׮�{���r���"��	F7��q�W�8q�	�h�yd��y��.�$z�X[?��z,�#�S��_~4~�'^g&�Xt7���%�4����Z1�Ede��u�1X��'=����o}^\|N����
��]�����4�����o|c�Ź1[c�Fg)iتШ����LTp?M�u����>��kC�a�C��*�Ep��V����g7�q����l
i�LJ�7æ�0����7���QA��@ 0����̉�#�٭���WV��a����Kgq�<՞Ĥ�FSWdXAn����>Å�o]�O�l�8��5������(0�gH��0�Y��=D��'Sd^^�|'.~M����6��_��ϻ�D����쫊���|B�N� <&�(`.�*�,��:��TIhR��rEG���f0[l��j7��ȶI������X��2>c�(E��9��er�~�S�aQzȜ��Nk|r�69�i�gTl|E�B�gt�ވ���7���[h�=�ɫ�:��"�r`��9[D�'�0rKK9՟1��y����L��{�f�������j��T9KЋ��"�/�ѡ��;lU�zF��{�$Xզ�N�<���P��w[{	q�P��})�N���jJ_�|U`��F������
�*�-}.ҿ�_�ò5�����
��ן��Q�T�׬U�
|�W����3GA�C�5�'�f�χ{�Mu9�~�r~�<��A���.n��{%BaO���éi,t&��R���p-���\U�m;�/+�f������Cۑ.<ύ�_��R�){��'�L�u�*;�8�͠�{��֒sB�9��"h� �	����7�>HSqAk�V
�b�<����=
X�J@$��	h�ؒT���Fb�O&�K'e/k��F����������|{;��љdo�"V	�G�][��h�$5����L�TY=�]��B)+��< �]� ���)�� N	��Cr*�"��;�'���x)y���gͬ����)��_W�������j�A'ӟyS���S��ǲۋ�6%�Es<�Fw���nxF|�C��p�\��Ićo�3>�[�{�
p����a�]�_���\g��i�[�u_�����tK�wOEg��x�ï�����������/f�}z'&�DQ�"�n^�M_�%�D�Q�>�3$�Y�f��cZR'���At��L&'Ӝ��5�^{yZ#Y�S�c��  �sUГL���s������up5>��ؓ,�1�M�M^t�H�p�bB!cJW�Щ�̕q����y�[G��������p��V�Ґz���3��ُM��h:0&�5Wb
xMF�,U43*Ӑ�s�D������J���fbz@�D0�6��p�J��1�t�/�{{�����8��/r$��F=	r��"�� �X�rvV���Al�������%����$��h�2�î���o������������E�t�U�
��bb��խ@��6`6)�Q*��Z)���a.P�mHx��}�>��A3?`���5����go�,g��8Z_�����F�F�8fR�#WX�E�i~.;=8i�:
��yDp�H�T����W ���j��*�����_���ޫ��g^�@0yh�uu<:�0�t���j��Em����Z1R�Yo腑R�3�/F���P����ٶ�����4"Ψؚ���{�qXtxU�7ޣ%�F��2�kq�DA�ō؃� K ��	h�;m�����v����^�ǐJ܍��l��e$���`�^`�8T�{k*��ԫ�Pw���Z�j�΂Ǣ�[�H���qb��h����Z�����>0�cY[=����������"���ό kz���>C��uk�r`�7�>1Q���8)�2I�=�`LA5��W{��u�:���B+��R�����.Hĥ򫪉�I�Σ 1�38��OL�-�&h&Qm��������k�Ne_
0#D{��I ������
!3��!�˨I �s����eO��_Z'Y%�,g�&�8+~�Cɗn|G11M�΀S���B+�x���w�1e*Z3^$�mr$��)0�J.� �|6+I�,jt#����zY��m����k�ϫV-�/���;!`���@�?��*#ZN]��J*����m�������	�:� ����a�u�מ���?N�@��������8?��gx[�T�ȗ���d�f��A��;���g"�4��t���Pgom-b0��r�|���bS⼗���d0��}	�39%P�I�n�$��QVK�OV!m�_�5� Sڎ�������x�_p���/�������b�[D�ȫ~5�y��%1-_ه89��b?�ӓ��_�9�_��q���XB�I:�%��Z�M#N��O��g�?�o[��˽���}��_�9��^����ŚęSgb:��́��5�/MO��P�ڕN����|
E�T�d���%�x5�0�ݒ�Lf���su�:�ְ�R(����Z�tP���[���6�{}�{4�Y�g�Z���-8�)��#f�=�]�0�X�Q��Ո���@(`�P)�����<����H��"+��p�ϊWJ�T�hM��|o!�i ��Gz�AVN��:e��w���{/(��}\p~\x�8����bm�H���?�^/���[�G��ĩE��H���:1�g����/��^�3������O�����S���I���������v��G~>vGc� 1��&P�������-	n(�Q�9�ˠ.�\��Ѥ�ڛ�`�҃�0��&�S��d¢�4+�NL9��aL��fR�~�h��X� <a�#���,����Q%"� p�B���1%7�a���SE/�P�T�v��1.��ڀ'Yg�Ax&�H��J��x�ױ@�)5�B7-��}���>����'u�
b�N�p�����	�,`�L���k���H��;$tU=#y��%�/t>&����
�SS7EmrEseS�Wz ���I�{oEW�i��0���|1T �>��30���!(A�:���5�@����
�)�b�0_ε'D���Q಩
JZKEѠh�N ,`{�h���?W*��mjhur�"��i���P*Y��l���� �v(9D�p�������!�V������m%�ICV'Y��m���d��
�ro�D$��2�1���9ܛj�%&'���ZxG�Je�����R���W<���m}��NV��y������z[�.���=��"kܞ�7� ��"8_:C-C���ʝ'��TeZr_����t�K��"'�4+� ��Z 2�7	Z��黜�4UPh&=���)�T������jV��|�g��s>G����yjڰ�ճ��.D�6�{C���	>C�.��~�ǆ	)}g���$�k��`O3�Bjm����oP��H�F���
H���s��yę�H�M�b)��>�*V�4b�`w\�U��4g}��� ��w�X�ro˝�X��Dg:�n�"�f>�F7箏�b���4�[���K�W�I�qƵ?����ӌ�0�ݭL-��.���	�3��d��� e��z��8؋������q�������u��z*oVL""ŏ��k�K�����c��P��<FY]�f��,V�19}"ֻ�x��O�S�+/��� ���$M��ٳ5����A�tۧ���#>z��&�    IDAT'㦛>'�?��,:��.O�3�����o}~\v�fjj�	x��N̦ԟ�A�C���kj��l����UӚ��Soǿ
n��A���o'�~��u�
���E~�هci0�1{|f��Q6r�t"�����E�Ld��CV�M��$v�#2��~�g��~���ရ��(p�j���+�y�r)4� �!Jn�utf��@Ƅ\��p"_�\yurd0@��<��	�ԝw�]��+N�>����/��.>��~d3�����b|�؋~��?��_�3�X�R�w��n7{RU�*4B�Y,&����^O��~2yGi?���n�0f�x�O�������_C�!e����ŷ��k��t=f��>���p�M�<�'�a����d7R
$���A�v��0z�<�CRe����Ys�g�.�*)f�Ru7lJ�����K�a}=����Ǳ�
[�����iV�dK�X�j�j(�~���t�	�4w�8�L$\�Sٕ�LI��$�	�o+��V�Eҕk��YPP���J��)�PА�W�NU#��R���"G=]�S�݀W�I� ���cد⌅�W[��
 @r ��н�I�r/ki�Tx�,�[R�z�%i�R}�}7��@�-�%���	��K�� ��m*x�H�:+����2]YU�<U�ƀ\����Y��]��3
�UG}9�d�ƨ�-���&�s(	h4S4k���)��Š)U�Ze���I#�|R����h�A�#��V��A��ζr�T���o��I^g��{���Z�+�
�UH��Zx��*_��,<�����h׽�&ZgЖ�'�;Nh�`�����m%��@����0�n[t�}}�L}�P!D�z�k�>`R�4O�g�cVt�h�p� ��F����2�R;͂iž�=���gbQ�m�	�3��	���΀�@�s�_\v��A�<S��+����5�/+S�y�8r�,�j��1�^H&(���4�?W+���H��\4���U+�,���l
��� ��u��@[��r�b�1n�H�0�I�ׄ��\�l%�> �T�D���%._��|-Wl��ǻ�oNJB��TS�r�MN='8�*�Z���	�,�kD�' ��Vz���<�.��B�0�[�!�˕��$��D�M|b�⫹&[�V�I�� �{HN�VD�R�%����c5��<��LL�s뵨��Ud����,[L&�7j�R���e%0�=�,Y�ypd���P����)�!����$�[�;8����ϋk����sL��&��G_�_�c�4/L*T��Ǳ�N��/��N�b�Tt��k�|صqds36�Gc>M��^<�����>(�k����������x럿?v�V�����f;�b'�:;��g<9^����9Gc9���~�9��ף4�:�C����i��Vx� �c�)āA�����:.fQ�Dω���6:�&χ�kQ`���Q�%�r[��hd��2c��Jȩ��6D4]2h��:�Τ���9�IU�=Ɋi��/:1=�d�
V��;�l�6�G	)zf�t���*W���6������^#�WP�����*�+��d�d�sa��i8wV�2yZ����T|��Oę�g��^q�eq�%��%���t������~���M��������w)��Hz.�9d��b��~�V;��ߍo�ƯFb�L&�N7t����ߟ��3"n�?�E/el!1���L��wVL�C����A���jHU�K�lV����G<ꠧT��w�*��ڗ���jJ=���ğbG
���Ytb8�F¬�xK,}�y����He��L�q���"�R�Ya'<ˠO� WX9!�.�^��fU�J����R[��ݖ��d�H	�H2�c�C�Xt����+Qv�i4�I(#��g%��@����0l�78nyg���|U�j��v&��|���򁉋vg�>������*���dX��hz~�=�AlM���91uo�n�����*��� �"��̕A��P�v�;�`�M���}�Me{]�`'涩�B?�<�d��[z y��-M��C�{�$�qmc�2p��+�tb�u���GvE�I��jr�d;����T*�$2)pVsԐO%6�Y�z�s��,�U�=\�7Z���(��_:/y��v����{�1P�0��Z��g��o��)��*l&�>��0�〚/l���ů7�dJ>��:�Az���(�����`���)Y*���p%gNc�ӣyl���%�����$�De��h"��;8^
��#[�TZ-&~��U��ʼ���y��0��O��z�K�d_%��=@t`�Ԟ�6����!5vIw��[�4������T������g�g�f�S-\�7`���r���꽪���jaKP��"Gף-JU`z ΉM�+N������@FӺeh 6ǳk͒��mZ�@�*�.�_�.��۽�
HkC2��I�@T����Y��<��(n�g���i�ډ�؉�"���r�It�0����}�:���r�Ϙ�lDg��d����c�-zS]=&�J�9�El���3�Z�4n�j�'�9�j��8~�^�U�=���='�����A��NG��L|�C�#1}����>1��QRy��k~-�~�*�:8���t���ӱ�uo�w&���G�_�yq���w���'����� ���'�W}�����n�|Ս?{��������>�=���Gb-��|;ֻ���g}e|��Gr�c̩Ȼ�I�+󣬺�AP�%W'�5���  ABs9L��s��7�`E��A̟u�:)l9�ųI+m�s�= e�4��	YC��CȠ��=P�s��.�+��0Ճ�M��D�Ż�X+�I�k���Ŋi���أM�럅�uAn�0��8bvR��&�D�TP�|8TUHݠR��;�w��]B$h�%I�W�*��p��L~�q�m�[o�=v�w`�����K/�#�6c3�yG92&/�Z���������ݵ#�c��@Hz�F
t2�Yt#����#��x�s�2���~i�2i)i�ߐ���|�p��`�O��x�K:�&��bQ�4v�	��ڲ�tʠX'( ʉ�H�H�r&,g�RX�0M=���y���UJɟO&9J��B7��� �Y?ʞ��2��U�(M���ɴ	�0�o5��H^�'�h�L�Kb� �#��"D�C2=�-�CfBk7|��W��US��S�E�X�&n����W8CJ���>�k�`3J�\���/��� �������+��B�7�@����N*V�9���"�;9i�00��{������Ē��Q����	*��D���P�?��R��x~v)FX(�23�B�#pǈ�=s�� v@]~WB�$�'���A�Z1T� ��������Je��Õ�ZR�֒I`����WT�fOb���~+�ՙ�pY�S��;)�Jq��h�Y���O5t�U�ĢO�#���^Qީ��<N�����dW_�s��j�TŢ��.�J��`���ZJ�+�O�U�D���LNywH���;�'�+W0U���a?_u��ӡ~�J���{zO�$3z☸ZEuR�+�d� �T���~Z�P]� �-#�eZھr-��z�C O	�v_V����v�:O�σX����Rś����8r�$��Gd��	�m�A�]�m$����f����q�� �i��u,2��TM�J��;�>�^���N#@T�U��1�d�=�X�Ӹ�F{�	|���(��
6��E��E��l�u��:%�y�	L�]�g��[ӿy`l�u�U�4;�UO��\��|k�ˌ3�D����F@�1���'#��<[R�&D�뒱Π3�a��|��A�"&S(���o��f��Ie����e�R����Jō�7�lP�>H�4Gg��b�,:���%Ek�:�:��S*��c�h
��6�\��d?fۧb0ۉ�^}a��{�1�mӪ>�ST��ܿ�����7�m7�{���(��M�M����Әm?O��ώW|�7�edi7⎻���?��q��}��_��x�W=!.>F��oo���D��}k�៾3�wRy��n�b+���_���g�Z7�f1�Lbw� �$��Nt	a7:���hR����Q��L��I��TkaL�\i�'�s�pEű����5O�>1g���T��(�QmNFcm8;�|+�O5�|��?������]"M�9�u�@����i[�9�|����2u�Q�j��4R�ˊ�_�TID� �� ����#�R������R0Q���,Qi�B*PM��ł�2�[>v[�z�m�aNe��.�4.��xlو����3��1]�mu{����z|���1ؼ(V�DO�1��|;1��c�u�G����gb�����'����H���(/;���O����O*��E���7��t#�a̗I�M��'��A��HL���sl��:zK�U!te�w�T�t��E	�ݤ��`�A��Biމ���{1\K����E\u@��qAIWcՇF��$��T!M���d��4ϙ�Y��L2V�A%�T�x��M���s�L�������J(+��S�����U�R*e.���K"�s�ڔ*#@�O(P��5�B�̄���0kU0��P�9������t�/³�"����iI�SIa��%�@����%��;Xa�R�u�ǤWD���[-Qa��Zx��gs�\u�(#S�T�g�)@S�ȉi%0Fk�������\��L\+�a��II���H-��	P�~� �>&J�ڞ3-\kB�����O>��N�E���I*a�ӭ���`d^a}	4��v�"�U�^�5�Bk *�s�e���޳:x��`���{�lBk_�lT@�,i���!��P�;���#�a�;�>��^V�<��3��zy�@(	c	�'�5�B�4Lkm�b=$~m��D�����گ�MSC"覵:�JG]n-n��3vl��Q�6'�\�:�D� r���l\��%ǖ���V��\u�w��Ň��
�X����]�%D�ߴ�K�@B׫���v�G���k vr�.�gN-���n� �0�#![e�J�*ﮔ��(�V��>�� P�e)�]xǄ3b�mlb�`�
h�g�U*�ECv�D�kh��r� p�WE-Ë�����%�Ctj� �o�۴}�G�)�3�2+/�шB�2�I�Y�mY�H��Q��]��.;1Nv^
 M�1�݋��[�hϜ%[)s�P&�y~RP�JÊ����h	����9��ޗ�N�C�`���G�[Y\���eX;�ߓ��~E����=$��əx�C�#1���ᡊi�c�JL���f��fRy��P!��Nb����Ĺ�y|��.��%�u��#N�E�ȿzC9r4���O��>�D^H���Yćn�/~�W����2)x��c�ڊo{���nxv��f���czp;;�p���#�*���H�P��#�!�*�Uyg�`h���<�2����R8(/���wՎ�89/�8�DR|l�j�%P,��<�S?�F4Zl��y7��+1"q���z}$��+�X-�?|Jӥ�<���C����M_=䑄�ؼ"��7V+���5J�$#`$�mzw�(_/��6���1�����ܽ��h��ӛo��rO�;�ܸ���q���<L*�hǱ?�;>xG��7�F|��g��ya,{C�F���"����#�����,����/���_��m7<-�݀Y1֍C���G ��ķݽ�o��W��t��|�JpY�y���#���D������Z�3	�{<�#qD�@B{�|��B�͊i��bR�}�9_����݅Q�e����1��uV}�H�D�_�
B���|�t�yw�=&3$�@'Å{'�:� ����R�J����ǽ�xֵ��X�Y�*&�XL{ԬB� vBQώ�s&�sִ��C�פ%f�G��01��l7���Ff) �ȩL��E$\�n����/Y%bb����2��o�լd�]�ᒀ�޵��=�0�͒�%�ЈO��5!J��:`�XvlEp"]�3�M�lG3� 砰����7/�I���[%g����>iDN�\ךX�N���`R`}�T2�[�X����Z�5U�]1�Y�}>�hj���6�3����A��A���?FJ�J$
i��WZ�xhU�J��ERy�_%����0���&`I��󙊠���x4�?(Q!�)���
U
�>�KbZB\�T^�lj��X��;��5���U������ؘ�颳��0&�V ���j�d������6�<��w�?W��Tmm�r-���GuG�K�Ψ��Np]�M�����������
 Y@ϾeLV|���Pa���徤�HP~A��Uc���K2X/������&z�k{�ʝud��;p�q�*��Z2
8j��iy�P�-�kR">��m�D%}�f8�ƞ�~����y�*$T�檞A�v�ۢ�K���`CR_G:�QdEB�*�7��Lb�(ֆ�q��������=w/��� �%��'3,�\��h�H�`�5�4ִӍA��U'��^��4��I�=؏Y�;Þ���[�j���g�
H!8b
��f���"K�JQ����3J;X�44B���nָ��ď���"�K0��ݭL��1W������uP���C��|�\�;??�&�;�"3�^����n���b�܏G=����}}|�UG`'����uk���O~��?z�#b3uL<�G@O.��$�w����?�8u��l����N|�?yf��%ύ�~�	2�흽B�`մ����F������=&�hzg2P� *GyL�����*�ym3�mSTSѧ�.aML�A���P�'�P��j��@�(3Y�;j��|q�u�6F�ӡd�(PqЌ��s�J�Fȳz줴Mu]�tNgxvbZ�x%JS�hu�V*Y��9PʿfЛ��N���*&�-��ƤI�V���29��`�ǎ��YO���⦏~N���_qi\x�T��d���Ggt,>���U?��xׇ����X&}w0�A$���R�2��1�Dgz2����������=\DIg��x�g@����*⣟�Ʒ�k��l#��	�����i)=c��ˑ2)s�=1�g�?�|���� pd�+e@�^R�K��F#���o�>+������ps#����i(!�!��3������	�|	���4砲��Ҡ����� c0!m��<�p��;�����Ҡ��^�d�$&Pz�h׌�#A�9x(�� ��v�K\K�y�,p�U���WIzP�ֽU�w����qS`�A��p:�
lQ	�P���d�Q\��ߢ6J�*aW@��c��X����i���#Ӆ�~\31%�T7�sm|�lG��gȄ��f1�ZYk>�qT��Ш+��{�~6*�%_�FɆY5�Lez0�[�?W\p&$��WT�d��D�Ac+��Ϫ��$��M),U^2JO��+���������7�WM2����`�A[���	�����"U?o�<<��@-VsܯT�u�}��;b�<� f������5"L�;�P�K`k@Z��U{�˜�h��^�$R����<�9�u�\w״@�y��$9d 9r\��N|u�l�|�+�Z�����6���"$�
�[����#XA BN��Fa�QF$�Q� J����ۭ��3ʻ`fEK�|�9����;S�d\�Sa	V"�@Z�?��զ77s3�0x�W�1g�>#A���m�jlwq0?�1MS 0�k���@Jh
�F������pf��6����i��>��������Q�i�l9#���G%r��٭��X�<�hUk��f+j�RI��{U�.�1G��X�"<y���` ��38%ޣ�2_�j��C\t><�I�>�d���H`Lϋ���}sH1Pg4�#F�&֥���w[� �qx��/39�b�L?�o:���>�x0z(�k��At�9r/j��R-�ހ�.
1	&>��qU��#�!3�P`����G��8 :X9e���g�݊�l7��c���~^<��Sj>-1�F'�_E��k���{b'֐qOg3$2��f�pv&�����{^�������F����� &@ٿ�qW|�K�I<�s.�����5(    IDAT�8q��x���E�r��ꎃx���P|��O�|;�:g�y�xr��;n�s��M"G�LAs"�F��\8��ǳ��e_�)@���g���eJ\�~r��*�)r0�~T�kt���m���J�5j	�yf�y*Ȓ�LH��X���;.�� h�LU�=aD�d�MJ ��MAB��LL�,[�T5:���g�U�,[MN��S����"6b�)ǩ�����S�r-Jx5A1
٢e�<^���R��?��8HN�|�;?�=����މw��q�m����8����+.Ei�k��b�ˢ���ޝn��k~)���>1<����T��>T��i�I���*�2�Db:���T<�����qC<���#A-h��������9D� ��m����bwq,ݤ4�;�7T����i�3pK
�h�>�D�����H`Cπ��L����Py���O$�S���`/���x��LJף�2�� t�?��� �U��/;>���?���cn�,�Y=U�&��q2FPG�ƴ1�H�}/���eR,�g7@�-�N踪���-e�7�٣8V�o���BW�*ּo�x��LJh��� �25<��o�(	�����0�w������E�������¬�� �;�9�t��� ʥ��l�ޑ�؇(M-�:)���昙ښ�\��~��b�j`��בy��$M��V@@�!��̽�d���|.U����!`��PE�E, ��Ķ硱�`6��T��Lz>�Gр����
��q��0�Gk��U]h���y3K��X��'���X�l�S��L%R�]��Ժ�W
@u��SP"%lP�TE*�Y\�3}�hNnn��Z=R��K�R[���3��(�&��@W�Leܖ���h� ����Wf�UT�	��U=&�bob��x�� �̞>�ݘ���9�* 3V�� ;G�.T{���V"�XL�u�>8���$ep��U��s6%�A{(���_EP#�h߷Ġ��ٛ�)����~�ySw���,;���P�ENN6
j�Vc��m�A#'f�P�_/U;�5Ҽ�=(X0Owk�+�
fr�la��H2BQ�<�;�>h}�C>��u���0��p� b��ś�A��{�QlI������h��R��)�d@v T�����&�X������&��JT15hQ*���H1��R'�����W=�$0�q������X��xF�L�����d0e�4��lo?�{��M����Sr�L�]���S���0���Ҵ�Ic�ū����G{o�jV,��TM�1��簗�څ��l�T����W}��ǉ�b�Ze=���u�5��w�v��FSl\J���p�_�ŏ����̸�(������_��8~��x��W_�[��5?��[n�'|���s���8��R�ݸ��2��~"����c���թ��/������0.��h,�������ZTԉ��
=O�B'�#Y+/v��"��K�NL���D9]U�u��q�<�����j��ʣd�b.g׃L�őP����rf5�AK|�cc��j�)�^+�nj��iɦ��Ǵ��9�|r!amRJGS�Nx�mkρU|�`l�興%ų$�rb��YY����)cNU���Ux�k�3ɼ���n^�
�{{H"�_tIlll�=���|�;��=w��� 1����1Z�e�N�N��������g%~�O?���KlD���ɬfR��?w��^'��Y$��=�a�ĕ�e�����ϺR�L�'��w6P#?���T�����_���y��\�Xu����af_�)f���琨Y�_�b8@��%p�g�}?F�ᴒ��[:��bg�p���&T���F7{U�S���0%)U��^=��Ms����$��'���b���6���h�.{ ��g�t4p�{E���g��M��ji�h&~	N幒N��%�E|Z:|����+q*4�k����Y�� =Wv܃��3ZU�r�������#V�-"������'V:k�ɨX4(%y[��LN�{��w�0�b�e�R��Kr��l�>e����Nqk��ek�/�V�\#&f����OÄ�(2��,a��VK}�AE5�U��� �1��Z�r+�00�w�	��ͤ��i=גWY�H3��k�Zۢ��P�E��a���� | 0&y�G�A��աI��7N|�O�l*��Lc�))Nz}�X>��'e2.4�����I�����<�z�P��̀��&���E�Դ'H���<�J|q�EkS�Q��3�d:�+M'Ώ��> G�a��@��&���N����|3A�$�X��*��D��yn��@BbP�������3-`�WI�
�E3��C@�A.W��I��y4L;��g;�ǠA��iDCKc�+�k�� �}v�k�������R�>��x���<&��5GE��q�L�8��Y���x���A���i̚F�4=��3���>G��Q&r����: ��WT�q*�У��X�ad�bi,�5mr*LD<�x@ ����0@E��:�8�;���(ı5���s"%_υ�T�Z� Л�ɤ�ˮP��p�Y�>�`���e��@��5�e��EJ �z �c0s�s��l�Qvy~����d<��1�"��!'@E�)n��3��>�|ϵLޓ�[>��tw����2��{��H�Q�=TgQ0�Yඟ����b�i[礃)�LRK�v~M"NPV�1��$� ��ޛOI�m�g_��~SSy?M�(�I�l#�'_�����"�c-��^̅j�3X�ۍ��T|�>+�놧ǃ�qc>tۉ����K��G?:��+�4և��Ǐ����ɻ�'?���9O��X�-Пw�}�x��D|�C���n����}m��w�(��+b��`>bz0��!�h�������Z^�(�3,�Ã�'��ʄ�A���#��t�a*�A#pK����^� �U�.qG*=%/�U��hnc&j��@l\]ڋ**?��z���<�?ͯy6�pH�l^МI+USVK5��PŴưx5��P� pReC��t��,d��#�Y��9������#d��&�IO����C߱hx�Z1��f%�ywgŰc���i��x��{�q�E��ᏸ>�=���d�m��!�0��H�0���w�����*��Fm�*@�r��q4NQ��$�IL��Y�W;q��,^��g�?��G��T5�����4���^�gA�;1M��<�U�{K��|0�XD7uǱDo��-���OJM�a��YC�'h+����9(�>���D1)+L1��Y��Ĕs��(���Q)�_�S�B�qW	��P������w15��T�M�I��Q�0�7�G<���Z��؃��:��w�W;rVk�
�ĔI���FpK��8oh�Bd�iJH2=O�C!�t�N��[5?N�a`u �3�]a�H���lh6��j���qϢ��1�2͞��m �Dsr|�J*���S��:��#��4�%!|[(�^z-]%S/^�Z EU��$':�F�f$�����	:���(ބ��&�7x��V�Uȴ��0���Wa)fJ��?�`BU�W��#��m���ہy[e=<�TC�-�L��,-��[`%�Wj<�
�dZ��SuKG>E�2*Y�3AG�+Iv,L�#�-D���[k��Xi3�O喥J�^?���sù�P@\^,���7��AurEA>;9 1��b殪�x��ę-^��Zz�H��=�N�<S�o���(���4��ࠓ{֋3�����,�ҧ��T�jh�g�
u�Oj��u�\Y�!�#vi$�}��E��R�י��Ȥ����OU���8�"b�I�W\���hPN	恒"_��IEƒy���+���ύ������������^J9}��Cl� +��@U=8�h�	)9�x���Uh��6<��u=�͸>Tڴ�NB���>\�:�,?�<%|e-J�I��\?���DU���d�����Ƭ0�����ַl2�jk��tNXk�) �l�_�Mr�I|	�Y�Jm��/���&S��88�xbGl$ ��Skm�q}��L�3yԽ=��Sc����.�l=ZNb������ ���� ��*���v;`�%���ee�a�~��c��B1Q�S����?e#C�w`�$�Gg7�4'�`\�l;>�ҍx�+�;>�qC���G�U��N�"~��o�?��Oƙ�8��'�)�y>�Ι/���+�O�>����e�z���K.��[�a:3����}g|��;�iO��x��b�<�Ủ���U��|"V������]v4���n�/��GǪ��E�Y01M:�a,zK=4�2gp()�`*�S$dLLٳ��QoiP��2y�˂$v��LRBS���a6_�L(�0����a6e
��9+��&�rϔ��	E���(+�5���mmEF@I@0�߇*��e���i�"UOeC�J'���,U��*Ez�~R��w`bJ�/��\s'����?q`嵴�1w1�����>-S�9boo�ݍ#��^G�n�y���w��n�9��^\z�Eq͵�#ǎĪ�AE,�,{a.g3��Zŏ��������Zt��'�5�h9"�7�="�zI	��l~��4�݃8:�ĳ��K���$�Eʻ�':B�+��������LJ��:�Y:�n7n�{��'~.>v�<����KbJ��IКL���z&�kl�o����J=�@�ݘ7�$Z�Ӳ�J�(%@�*҃�M�1+�	��K*��P[���'#�� Ѥq�`�`8�v�
�xkG6c��*¢�"�
�
�ZS�C%Z� E�Pe�爁 ��3��{�z�+;!QS�P��g0�Ab`;S�mP�d�������g,I�2-߂%�V���֏���,^T2��XDI`a��>栘w!�2�ސ>�2�7Փ�d���2U{r�!ܠ����K@�d�UX�[
�����v^wD�?�6rE%�I.�?���'�&A%1��4.*�\rE}ͽ��b�p�ME��ݧ�퉫I�d������U֊���`K�n�ĖqU����A�U�$��re6=�lQB��)o>-΅�S�Ȓ`R����IK�V��WQ�qh��϶�Һ��q�V"$��eb�Q�GF.A��V�-�*$�ςKT�6��z���r��8ö����아����$�R��(��P��UA�m��jU�}쾶x*@�FV5��tQ�]���>-Vk��*��I,4T[i�O�Fk�wu��>���3�Sb�̹t _s���>6P5O��*qJ��eb���l�E\w�5q�5W�����7��l8l@@ 8C��=�ډb�����3�=S�i����_��1]���W������~�m;�`��8^��1U\�Β����V#&>sƧbS�j���ؼ���AP&�ȫ�;U�-�m�����M^6	0{nm�h�.�v�E,�r�JA�A������2V��JU���Y��5�gڔ�Q�� bm�,r��	p��.N�M�D�_��a2O�݋��cr��0:�^���b���S3�ԋk��e A�>�+��܏�_gΐ�S:2�rR~����%45 :G[��4�*w���f��U��Q1����G�+�iVL���^�c �v�t���/w㳯<'��%�8{�q�aY�����s��O���}���_�E��?ʼ4�݈w�|?���&>�{#���߿;.�w���x�3�2��<P,gb8����&+�v;f��rv�6	!*n:瘢��%R�K��RWOss!~4�6
5%�:.,o�-��cRȦmT�8��U.����{�>���P=�Y�����#:�"!����6�D�S]��)�� ��(I{��6L
�z�������S�	�r�]���M,�O��ɤ���oh�(\#r%��# }@�9���c`2)M���.�#��%������c{k+.<�����+��+.��(Ux����0)y��1�ǟ���c7�>>u�$�PXS�B��Np���t��F����`��x�C���~���A��B��`�0���v��&���w|��n�j5_EL���Ʒ����?��ι1���a,�z��*����I-���хq�I���B5"��^�Et3	�eO)Ŏ(tD�L�O5���HQ �3��tN+�����������b��S�H�.��-黣� ���fE�AgRn�����4f�s�3��mr�U�%�`�@Z���uӛ���	/�s�Z��r�
�[h�t�������Q�XR�j�)�+�"�V*4���0~��mG�L&�W�VY�\�>�� ��8�6�l	E�{���\�$%I������W�џo�X��S}>V�U%Ց[�1X���C"Ԭ";p��d�	�m�?O[MdU�k�^6&5�,E,ӳ�"��k�倆I�D��X��{�}R(v���E��4]�H��(OR�N������b"9��Nh���ݕ�CT{ku�1yy�S�9�J�TMQ�����b{n���J* hƾ�x U:���4M,���bܔ?a�N�L�K�R����rˠ�M��C=�Н����io�p�Ej���`��͟�&����4�I�� '���>S�1���J���`��G`�>;���>3��U첉Z��=�l����g��@�c�����qhS�/�ĩtC
�<������#k ��qo��}��4�4p��7qϨ�d2�Ǫ"ʢV�~��"���B�� :ʹ֭�!��O��P�>��2VD�-�'걷fF4@�[%��Z�B�u���Q������<���J��x%��'���s��Z�*ʨ�KU$N(�+b뀶�,V&�Y�E7���Y J튜2���������j܋��8V9�n�C�2��b���L����
ש֛wr��8iW'�ù�Dx�͙:��b���:{\�ɼ�9�V��J*�ԠrH�#A�LN!��51e%Y F��l�����_��]�g�s��u�F�����?��������T��ZL�w次�1�힎��L���3����|B\yёzcV�w#�����{�_�}��q���Ӿ�K��+.�ݽE�{j��7�|�coo��At��c��x���E��7<+�9g-&���f5U%;�Āj ��Ĕ�ZMZ=���j�m�sq� ������.c��%�Ө/gUф¯d�)���SU6�\��1��3��b#hY�	/+QP
����jPQ_V����	���P�
�n�Y>�%[�R���{.���]�}�Ҩzr�02B�����wrnt�k�&�6�ʁ�gy���������ǏǱ��'�v6�����x����K/���8��EJBr$��U'���:����?�����d�?�Ja����ɤc�Mh|��H'-r��"�λ9�Ʊ�4��%__��1j	t�B�8�e߆S{v;v�ܓ6'L�����"n|���%�V1�Gw���Ҕ����<�4:�j��ǡ�9$���F�h��P��|��)E%��pI�B��٫������X��T�����Imş����|����v��](�%I����k�n$u{�<fR�PQ%��4{^A=�A�� J��ym��fB� 
w��Aa��Z!{��zM��=t�^�B%a���,e{Ա�@ʨ�3;z|M��b�+H6%
Ic2:J_�P#ؾ���\�s���"Rٓ�>s��/Y�(�9) EIM6[�He���ЦW��@���L��M���ܺ��IF���~P�"=̘�"	��rR����yLy.�����9V�x�i6X;
p��/��$��4��[�,�j(p-\ i�9��Z|(g��I����yȁM�~*�j�L,G�m@V�J£s��P)�H@�ޟ��C�I}��k���>�{��-&�܉��T���~��~v0�h��g�|ݣד�cM�@0�K�:����*��k0�0CߣDʯ���zVt����@S�Nbf�iO�$_�ڞ횜:���5k^��~>�a�����sשh�%p��O�$��9y�������s��q,w\���{�+s�?�,��
���v5
ɢb�)癘^v����|V�mⶏ��@�    IDAT��y�c:�s9h [�@#>�����m �-�u����9���b
,Xh;���/2� ��;;f̷0�����N 	b$���k�v^|ƹ�{6l�<fM��``�^�b�Ujd".!/��2�4'�C���{��J&���8����f�ǟZ�t�1�t14�t��Oc�?ar��9`Y-b5�Fwm���.�/ю������0�� {��JӓJ�9�to`;�g5��p�U��xVY���Ӈ������r��s,�u<;�=�`9!;��z*"cL� $�{��3يG^�����aǇ��i�g21��ߏ?x�'��r�ijkٷ�����V,vO�b��8o�Oy�c�)Oz||��WE� �D|���7����;O@}�s�ŵW_�sn�j;>y���?w|�HZV{w���T<�QW�K_��x�uW���6gr�JߔJ�HV�>���6�ߥṩ�8��Ù�{^��º_ʴ�5��f�\kgX)>�d�l'�A(
��
�~U4�k6P#�Nq��,j2{��
�&f�#���H
Ͽ*_B|�<]�+LLQ1�T�>iU�
y�K	�<ܽJ4�����:�9h��:�s��nގ�"�H
�}��gÈ���E��b�$����#q�����/ �!Q��3[����;n��G�ر�q���+|Ul�{NL.XV!����o�)n��7��w����?��	��iU%x�|�{/�̈ȁ�Dфp��pB�Ҳ�.����X�]���ʡW٥ekYZ*��,�H�PP�$�I�D�d&3ɉ2czӝo������� �Z�V�/޻����}�;{�}�9��v�;K20�9�fNٵ҆����-�c2\Ewy>��O������cA�lVL������]�A	������]�O��?�K�z����yY�!b�ݎ�h'�8Di��	�'z$Pq��	�߀��cS�)��9O,�H�K*��zi �q@�$Ӡ ��ێ��$:�a��.b��3�wY�K�V�܌���]��f���r}6=�G�i�pk�����;���d��Y����Q����9>�l����a��d���!��������A�,	���ͪ���Q`j���������Q��̿\�8���$����B� ����S�R]q�\�:ETW�if�2*ّV�+�+��d�Sz�j>g&��R�ϕכ��RL1�U��\�Tk/asy&�Pv�``g#7�2|-��l�[�RR�z\a٦R��L�l����D���J(3�?@cN�3��D�W�ӠYĔF;a���<P�h˘S
��XƊ���RP{D��e��{��d_��Lp��Xz%m���׮�癤�Re�#U ܛ��M��j%�+J�[z�2���G]e-K"{��!Vw5e�r����|�U,�#�]d�8W ��ܠ�{�H�*�c�pS��qg��J���OF��h?ЃVaI�eV������zǐ6�8��U�l{f����#��S(QNWgK�5�u���*`�rr�u��_� ُ[�H9��]X��0߼�~N�+���a�
��2Μ>_�e_[ۣ��]�{���8<\P�ՒG�p�Y`Q���P{Ƶ,L8/�xGN�ݑ̻��׳����Y�bj��-�x��I(oT����\���(W��n�*�����6*���{��Wsj���)�jH���Is�uL�j��7t-���xS�����M7�!�:\wP	�cypk�
E����-r��H��A���U��p�w�*>����0rH�qчjK�/Z0�b�.�R<�<�u��qzK��������?�[���h���Y��X�~�@��o;��%L7�]���9?�q�5G�6G+��1�0}�k�5�K��c�o�����8��P�W�1�Y�=1�/~���Wٓ�����{y�~߇��;�!��,c��;;Ǚ�?|yv����1��b��_����8�ۋ���������WG7PiҜ�X��� L9@z8��R�L8���L�	L�^EQ���U
@`�~G�����u:4����){�*ï��l)��n0@�%5<�@>�+{���3"���r��~%�-3j���+�\l0����@h���BI=@R����<�t������,��@c����@��\�ٳ�{�����s�DND ~)��}�DLg�����3 �g�ˈ�ZĹ{>��7�|:�k��6>�q��3�^KIL72\�k���4���;~�/�w~���n�c�n����\G���Q&8�IFd�.{��c<\��`Wo-�'~���7][��u�V���w�g��	*0��J���!u~?����q��+��c�F�G���A#�| L�ћ��mw{u4����N�ip"�8 ;��tGLc �P[۱u��~̑�!Ø��9�^�5���f����Y�+q G����!�x4��رۡ��*�<H�FA��XW,,�����0�R�^�S�k��Z�q���2�+����ĀW�{'�%),��<�s!���0�W��6'5�W¥d'�� i\bS���"C���
*�WzH��Z���w���,��I�X���3LI\% �I�����̭���5�IS%�V��۩}Jax��ɘ&����ƙ8�lF?���/�����j��=�z}*L؆*���%�uj���Oz����f�-���h�R�{���^4W�x]��[��D���DFp&-g��+K�_	Ly�8ٶ\0+.n�)2�\o6�R�s�*�J�+��GN�~�z^GR ����y���[U�6VJMҹ�LR��{���7�
2�Ą�"����k�\5A�{N�*��?�D&�VW��#e乃����x�Sv勠>G�)�i��p,0���`���L���|��3�+/ �\��� ������ف8��a��8�7� 7�	�'���\M��?�_s��ۼ�4�4d�n���K��A׭��;[-����ʯ|r������;�7f3�:����9�%^��5Z9������ʄ�䰢{��P��4R�<��2�#^�Ĩ�&6��=�s&h��E-T�!5�p�����d�x_x9k�����g�J�~K�Oô��<2I["	;�|��w�Q}^g�Z*��T�1���6�3���1w�'�N��=��r�z�c}0��!�R �������?����m����9�sFM1�������,�t�N��`\$����;�L�^).*qQ�~�m�� R!�%0e!���q�� ��5}�Y�|/��K���2���>�3�����t7"~�wo�?x�G(�-�\L(�(��|�|�t7F1�S�U<�+�$��˟7\s&�&۱�w��u�","��N�y������d��O^���8�V��46Ӈc�c�8�ӷ}<�Y�80#%����,��Y7 I�z*0i&ڼ�"]����dDL>�h,F{<�@�@uPy4YBz�d���ӭOQy�|jz�4�8,��Tu�YC��R��&mV����~���ZhVK!�� Y���KUOSRk�
��K��0%y,�T�)|^��dZ-�m�sr���)+a��æ��̓�����m�1s6��avt�최5�_ ��w�e��]��\7�����G���qx�'ƹ#q��x�;����Wƻ?p_�&�����X�[�&x�RB!�9{������FO�<�O6ѝ=O���ǿ��g���:�>���օ���2���f��ّE1�	N������b��/�0�y(b5�*�}0nC�$r|��>ݭ	?Hx4A�6����
`�^o������4��\�0��Y������p> �
��ɔ����ȵl��}!��ق&��^7F�v輋y�}Hw����q���LD�ʨ��n^����n��T���\'�	���B$QM�+Ye��լ:�*"�7���+&�
!�N���"�I�,�}|0g,*�W.O��V'�_H4=lے�|6�%U��m��Q������j�eɊE��Z���&��h��>)�AfxHB��' ����bv�d�-�p˧^У��8�0����JuQ��N�Kt���K�kI�%u�q�+����ؚgR� �=DI8dEU	b�6[��6���$2/��{9iS)�Į$����ɧ�[d,�~�
Ԝ� a2Ϩ��ә���Z�/����~w�
&�9Ӱ�����(�[)'tŇ�8	���^KNi�kR<��i��-	o�r}�6I�G(IV[)��j_� ��fŮ|��!�v��mʘ{�y��*����A���	����6���Պ�ʗ�+~]�+�lnd��e�I��m"�҈��6��rbdl��(	F��O6�UI�@�Ή�����F�k��J��]����|}'�un�6�4�EloO���=6��{����5��&o�
1��YlI^3�O亴�Q~޾��_�|�4�VW�82I$Vye�Խ����-5��4d0����OU5�~���$�
V�i+���֮q��rTu�s�
~U�`�3��/f^%'����/3K�[&�ո���gk^�&MY5f,��#�٦#��D��`:����X�h���Lb�A?zۓ�`�+��ON5�Q����f$ߑK�dHyTo�Re=ȧr�ڠ LQ9e���4.����W\��;�T�3.�*M��+�p��Ir{��mg�qx!�p�$~�G���vH`�	Gu�9�R�_��7�+��a���9\S��Y-b�w96��,���N/��O�oy�S�Q��>Sb�|�U��E\�E��C╯y[���wĥ�Et0�v5���B��r���Ƿ?��ſ���ӧ&����/cGN̼��ɇPe�$���S"�O@ZgOl�)���(�Ԙ�F�&���`���	i�SN�J �)q0/	�5�-������t����H38,?prT6��z ��d��-����]� s���٬ܬ�Z�L��>ޚ����V5�yHJ4�7�1EcV��Up#�P�C��*k�Ʌ�(6��+����Y�����׍W]��>wO�?��{�w��-q��������{��ؙ�4�A�Y��~�q�}��_{��ַ�?���`5�����OD`�a%��Ƕ§l��$p�e��nb��ư���r7N�g���}�͜iZ'H]�;��k2��7�kD�J�FE�;ݸ������>�͉X��#�-�2Q��������z�����QΚ�6��		T���	��C��2�@��ˠ��loGo8J	��D�|b=p}�v򍧀χ�b�E��� `���tȆ|2!I��97(Ulљ��@�+�������c�e���v���$���<�k�K	��,�љ�[�3���;T|�^ӳ���2�n�	?��w�'I�u'�����/�Ѧ��Ud=C%�Va��h�Mahy��?�=��S��4rOm�i�:N�K�ÑR�vVM�Z��E���K�'W�*�Z�$^kW@_�rZ�֖Ƃ�,W�3)ͺ���2k�F�s9�Ɗ��YƧ�9(7�:�3���H�2?Kuc�笪\� C���5���*H��ii\��A%�e�7�U~����@ۀ
�bdc-L�ym �����4��Y9�(�cH"��g�>E^�����k�40A�W�g�%1�ʢ�K��iM�S���1$���FAy>x�����擸�ɒC%&!JU��-H&�El(���5]H�g���g�����NQ����PDh=�@��K��z�͐8b�2U"�Z���h��^���u��
�݀X˿�y��_�`���u���e�I�Y*��-���qx0�9�[�9���y�llɖ����ۈ�K�-�?>M7�\�w��L�U���\�z�:�0��a�3�ˌ]>z�3�$���Y�����kĮ��Ζ�Q�QUV��Q1N�17o�k���Uޯ���)It�*'�$	�@MT6罉K��e�	�|ߩ���b��ŰӉZ��1����)�NyBⳀ,��5��bcG�7�p���E$�#�Qϑ{ܒ�<69J����s�N����P�-A�Xz�L{ҀU����DQ�4��5��b�nԶ<�W��^�1�������a����j��̣K)�o�����o�`\\�b��3TՉ�,f{�b���Փu|��y|��|u\w\.T�F �|�XG6E¿-6{ˈ��x8^x˛�/���XϺ���j�pl��c�8_���_~�w��=��c���Y��La5��
b����ZBL� ]� L�}��MQ1�LD=�� ǿG ��3u@7�/�OWI\l.��dypMNj�����[�w	���~����Q�=mÛ�/ˮ�z%�������N=.i�~L�Ur�ʭg��'[A5��Z���@��-��4����<�Q����-\�<�q�2��s�0��0�i��9�p�=u�t?y*��1�+�v ��mo}k����ƙ3g����o��p�C2�����e'n}����{q���s�;E��Fwx2F�c���	��	&��$���̨��ހ�	�'�t,�W�[\�<����c�puOcc>헏��������_;Z�P��ƽ0����<��_��x��^���8\�X-����I�It|�����W���L�ٸd>=Ȟ�Q��	9O�/�C���-0@O)�8bn�I��I�k_l�zQ-��FG��������t=���N���Y�EE
d�ԸGe~C)��UT]��;�/����CʉK�dk�V�f�4f9.#��V�հ�>+]Y���&��^�f&����+T^H9]�cp[*��&2�N�53�v��w�%]�)�L}G���=��±��5c������ʄg���B�q+�U1�K�B�7Ƞ�)�91VO{F.o����L
�j���s��*��u����M��ꢯ��2�}�$46q5�ħ�Nk�Ԋ�Ϊz.8����f+U��U���뉕��8zT�R�t��@����P֯$�\�& �`ϏPF�y���WV�э��)��-��7�+��E���TO������ #]/�9�2��©��K׈�n\��/d�%����FIe�X����f��(71G5do��t�г���z��)��l�DQ�ŉh�;�2q_/�A����K������H��|a��X5��˭Z7�ǼPr�:���Ui����Irm)�2��J��b^���E��[r�+��JmM���J_�cQ�D��fHzϐ���t���|�k}$[� �B�bIbp�c=��8�r�=����ؕ�I��#��R��ʵUj��mk��ã��Q���G�
�αZ�}v;�[ڔ+�I�k&k��Vyo��3���U~�r��3�9�R�z��~�rBW�te�{�yw�4fI��r��S!���P(}R��fK�۲\��q�#T�f��;���>��'N�.a���t[����T����	_��w��D�/(�ŬS�@#r+�R̩����/�t-'L({�{3s�TG�rgY/D��9��a�ا+�n؊����g]�T�R����q˭�˫q̗0���}6=`�tܙ������xf<�1�騄K>�m���˱�Y:9�sg{+v�'qΖ�n����,�%��x��so��ˠŗ�K��;����8>8��y�7�?�G�W�>M`:��|v�!�)¢��J�Q�A�	z76�1�ܸK��Z��|N2_�A'��HX��`�L��0���t�U�)�db�g"�m�<<NB�M�U�d*q��/Gld��wG�;��ecM`���5��]߫��3l�9+��)���N�.�4���=���<��t���9����e�Q쉒'`��*12#*6�mm�L����1_p\����q���1�L��/8�ƽ�X��M��d4��������>6z[�Jг�� ҏ��կyCLW���Oƫ^�q���� Rޝ�`~�dJ�˚���M�j�Z�vdQ�/���̣������������g|IL�,ԕ_z�5=m�迃?�*��1��'�@���a��n�@��%���\�z�1���G4*���fTL]�p ��*;�j�s%B�� F�`#[��(8gmξ�Q������=)i���éC�`���� ��|p��=~�y4��`2.C�7�PӜ$6T����:���s����瀃pVm��-��a΃���(Q�36@��W�!w�Ҋ-�1 1@ο���    IDAT��e]���{���ւ
q��f'<J�˯$���W�.%���J~�8�Ji[qN��	�b��j����<�MDJ
Fʢ^Z %���_��``.2?c
��[�8����,iJ~���}??M��}Pe�.sd�+����a�fE������QF�(N�7��aqޏ�WU{CU!�{xPʔ`$�� �����) ��K�G�.ձq�[f�jA#��:,�k鲜cx�%PHجZV���*M���� �m%��U/U��k�5q�7�/L��g�u���&�V *��Jm�O�"�����=Z�Z�O�녤r* �֪y }<)���Ni]��}I#'�pE'�Ĩ �HeGj����(��Bnd\0��*z�37q�v�G�$k0`�n�E�����*%	�A��\��u��SʃrZAΙf�C���>�GM>�u���V>U��{� ��$Λ��>K��caα�_AB��T�������[1����1���ݸ�8k�b����-��V3�E����8'���7Vj�g���32��Ô�V�����K����d%��y�)NC���'�B��������r�kIlbK�E{.�0��J���M�ȅ���kΐ=z�<o,1W+M*f2�P!['��$�k�<+:���ؓ�=��c�XG^�{�A��=��d4�.�t�Ʃ�2�y��G�=t���S8�.��O�Y�ZP9�{`�&( ���XU��!��b�
�t�e�O��4��y�6 �������;�)��B���W�y���K�Q,��X�1�vc����1X\��yң����?����3G۝E��o�[^���?Ӄ����UW_����������/�����&�Oߵ��g~3.<8�P�z?���������������q��ki$����jf�L�Uݡ���9N�׋�|F�] O�(SU��l�]ٯ�r8dՕĦ��ԋ��{,JBe��w\��d���b3�4U1NH�5���q�^8 ���r�"����̆��ҕe�,I$9�d�l'���ҩ�K��jE�
���:p8p�j��:j5����ܭ8K�Ńp����3��X�AF��9v"��wb�����D4c)c�r�}W��/o�z���������������=�G������hg�{T��z���9~����j�=���G���Ŀ�M�'K�Hl���x��l��lb��_��k�'������G1lG�UX��S���9
L}�� �N\>����<^��?���})b|:�Q�@���x~F6���r�Q��G��,�@'������i�şa�B9��81��`�Q)�3�΄���%��r�����BzUwD>|��2�)�,汜�r����M&1�ڎ�����@8j�:�Q�S�L",{y�8<p�	J��KxKS��{�9ƈ������H�	ʛ�.��qIR0+.l<ƞ��@U�LЬ��w���Q\��*� ��.�~W3�fj,cK�7�$���������?%�S<rE�`(�PK�]�&W6�b�Y��kۑ^�W")Y�boL�ƙ��`��@$Ly�)1Vb�2~ɤhv�fp��L��qRRY�>��'��䛽��� �It1�q�Eq��~]Ry��l�q�+��e�*U '�"P�����c����g���(W,��t-�,������Jc�t���*�-cos}J�Sz�9����zyƪ�W�@�LeϨU�Gٶ�@I-�I�5��
��k�L�`�s5��$\�	q>?^G:S�z�Ί�����+��{��49����ט�R1�DYGtU!8�,�{x��*{ �Ez2�'�K�,����Oʿ-����܋��"��N?�J���%�&����J�?�����!�f#(V��.�	�Y	�s����|VZHHDr�`[�{[���$�M28/m[lJdp�-"Ņ6��-r�/@���$ -�������`,�v7�[���L��gr����i]W��It�ײtu4����M��آז�>�b]��*W���6f���Љ�y��2�4#>	�3�iɾu�&�U��W�p� ��tR>̪�`B%##�nӱݽ�:us�~L:��t�ћ.bs0���.�/���e�������P 6�8wv�}�2��E?z�K��5������������p����Hn�Z�Rå�����j�zO�P9����_y\2ʙ��y���������~򷩘�7PC���W�����Q,�`���:�Ǭ�����3�������x4�{�8�<��S?���8�;��t�������(~���x�|_�8��N�[?8����#�ݻ���z���nl��I\����������ko�^�|��� ���u���>b<�f��%yCsV���^��d�hmL�'e��E�
U?�n����pE�,�L6��*9Aa���(	L�K�*�4�_13�I�G�d�˸5K*)���(� ���"%�bz2�U�h�B��I~�:��3j�k^�H����ϟw5���3e��NvXų�r(������#�f8SV�Y�x�C<s������s|�U<t�}q�{���A|��<&���b�s,�?(�'�U���|<��s��oxZ�=V�oy�{�?���p�C����D�TP��GU�	�|�^5����� Nwc����O�g�7Ĉ���"���o����P��GK�4���sep�:�vW���&>z�^,:ǣ3:�n�$U���~��0��?��j()/��ږ���}� p�P�<�/$�L�{�Xt64"�l4��yI)�A5=�~g/$��b�*:�e6�##����D4����8ȓ{�@����\J����]�yb��1x��3�3b�g�Ag�<��f����xO'B�\e�F˄��I:��pem��y��z��!���+~m�`g"���/ԂX�Ӫ�hnd>��+9�u�kaUN�	C�o�$�ċ����3��&��8���+*R�
V+8��B|i5M��_ő(�tJz�&���Θ�`����gUH�J���.{n�Tqؗ^+F��iz��Yю�}��EH�d�Vt��d"��83��3�'�F0����fOa�/�|�^j�zU�����$�
M;H��DFd*�*k5֫ɫ֘עi�p�%�늮�(�w�WZ��,S��������=�Y])=|)���)�m�;��hݨ�n���o�!��z��,x�N�9��6�\�_iT�Rgu�J�;�2�-g�ֽ���5�jN�VjWj��q\猽��ؗ@D���&	��[:]{��(�^a\b.��L�3�1As}�oքs#�����ze�H30c�n�&Xq!CI��I,�|N�����')g����E��|ӂ����'��%�31�h�����ވ�y�zf5��z��_��h�g[�		�5.�R��s����-�b	�ft��V��?{o�֮Bj֞fS�N�\�P�������^�y6Yj���gQ!53�i��X.O���)I��)��U)&ې���t�P������ὂ�j�`�+�!�n����#��U]����C���F�0��F�`��=�n��zQ���'��9�'��Y�	|�ӃX��5gj��2 @�c/��9��9�g�%�:��g�ާ	��^~m �	L��!���*�`˃�//`z�Y���+͏<.�w�����!�]�F�~HyL'�����{R��3��<�Dzo�������f���r
 9����N���<;���,F�~L;�xۇ�S?��x���讻�<����ѝ?;��x�3�)��?�q��i�n�"�C��J�!�Z��F�}�DtG��T)@�r�
���n�^�LY0\���!������))u��2�rx�1H��n�9�l�o.���ɔ;  $|�A�ϱ�R`Ƀ,%/%�+��H頃Ե>��P�B6@lW2�f<u��`y8�%Z��y�j�f���:$�I�*%���� ֣��?@_p_�{ ��K*�|��*QV��~܌�<�^Ņs���qG�c�Yqão��d[A8�0���H�΋n�����k��n�YD���?�K�5fG���
�
|U �V ���|��&���|S��v��q�d7���~k|��}7)yW���R��Wy#_3x()�{#3yʗ�jD�����jd��"��o�d<�_��B�{��38��@sH�)uT��q��Oe<�����J��V1 b�k�j�b� �ߒ�)]}�[#�w;�Q1NBbIym�n�6�GcHW֝�\�=`A����~,g��xT{�1>�M�.^{�<�弗}��5�|��i<G�z�!�x��ē �?�O�ku<��%@�s��f"I��5I�y/9N[鐦9Y%fY�>�w!R�"|j�:��*��;�	�ղL�|�6}W�psQ�Ӳ
Aֶ��h��+����)���Q�*�ǳ��/����]�z��S���J4�s ��,3�e�[#
	���̇t�ܻ�¬�v�ؔb:�J]Ju}�s�?�#�EtG�������oH���J�Mp��jԲ�kd(}G6Or��*�+2�f'� �cn�pO1* 0�ʪ��?� ��>��)����#nr�m���2�	��R�d��j�1%��׍{l�y���T& �$�W�WI��|��?���������s-{�K�&����</W�uW �v�H� �ґ&f�Vd��O���-��L��M�P�~���²n��W��ʸЀ?ʑM2xP��a>lW �Hnɡ���T]�}��~-�\�"s�f���e~���8@��λ5��ZQ��σ�xӳ�/��Y	ŢFWU�</<��1��U�M#��\?�A��h�?��u��}��G�1�������?��i����׼�\w��-<S���F�ƥ��U}�|���q6GU��TL�8�)Ԋcy��O �N,�Z�Hó�o��c���i������x/(%7�>,?��fb��Pz+�0+"��|��8�4�g��(�+V�?P����Ƽ4�r�	�0�%bp��bY���XL��d�1�b���	�Hw&#U6��^i)!�ɇ�#3��Q՜Mc5Üөb=�=�����x	F�>+��������쌱|�"�ٞ��S��@v��-�}�_\�'ް0?�k��r�P�/z�_�o��;��r��.
o`�4\���~�c⇞��qә^�����2^��?�;�;._|��C�^{M|��?!���>/�&#.�ˋ���~9~�?=7������rdLo�P\����W���-O��h��Rl1?�cŔ��d���@���	�b&�����C�p\.ث
i��p�xit��m�%��Ĝ�8$,*�"��5n ���*���y�jn��J�Q-t5�s�T���E��V��v�=H�)=���5��!=�`�I-}��O�Ybq�V�2���T<�v�R�H"�
��Kd��X���@P���tJ��2{
��l���ڃ�8�й��]w�x8�G��(�"�V:�T�0½;��C�W�I��Ʒ��������\E�`�;/�-~�W_������c��R�W�{VX��3)ҽt<d�L<d� f�c���}�U�Ϟ���UO~\�� �Ӧ�_5+��}��sU���%�XHe'A
&b�P%�H�{\ś�~G���o�{��� s�ވW*.U�0��U��칥.o#�i&��d��+�7N��0��#�oЏѱ���08b�V�� t�n^$�e�����`�>��R�١�e���$0nf�=V`ǌU�'�k��.� B@ρK���H�W�(�1(��1�LX�?��omm�x������YET�=�j�\SF�U.;n2�'$������>��l��I¥�L��ȸ�	Z������r�{z��H2�1��Ye]6#����8"��k���Vʑ�Y!l�GW�ZV<�a5Fy،����j{MR���+��L.5+�t��qq$i��j[��<����elguOϻ���D�-�ٯ�
z&��oW��﹁[�6��q�I�-y���{J�!s��4KpT%��!��m����?^z
K�c]o�d���Z՞L�鞙��ɛ-�t�����%��(��2!��@�?�AV��E�����U,�<F����̵Ǌl�[�HhA�?B��3�@�U��"�p�H�<�����g}����<�7�2S�«�\\u��f)���z��;r������K�p&���ȓ&��>Lx8���˓B?�1�o�nug�����>)�� ����I#����&�OK�0.b�f�lL��>]Uý����=W� >M����o4JD3�q�#�AN�j��� ���:
��>�%�$���8�gK���1�R�(���lZ��8B���d��=S��3��J���=�l��)�� �|0��-����7�{����sȧB��`O�VF"�l__ԫZR�kq����4{�Π9)o
����*?k��K�I
R�h3��06�A��X��;I+:����ȱJ,���1J�f����>s�R���� B��6=7�#���C�0]�	*���d���l?��
9RN@��!8E_��H��jƩ
��e�i��$��dR��`-�����_Ewq��EUL�Y30E(;�����w�������q��h��q<���s�>�Ͼf���+�����JRQL�L;Eh�YI�.E�����E/}m�{&�����>����8{�?�c?���/'����K���l?�t��U���G`���)�Ov8�R�S��+[V����!�(bZ��QjѲ�q���Φ�;���?g2�/��'�Z����O�j��y��6/q?C�_�4�WŇ�h	��e���� ��:_��r4��?��L-�ל��~�X�}�W49z���{>� �}�x\������J�dJ,��i7�n�s�}�җ�"�������8y|��k
`z���~������R^Ӝ��II��--M*�я'+2ذ#8E���
`7z�x�I|�?����i�����+y��Jn����Q̌��w?�I1tǡ���#������W��x��q��|d<A�>?��%$�w�(G���.�� h��b�Q����|I� F�p�e�6*��c���Q����(U��L��L���6=:��
��l�lJ��g�P��މ��6�4�� Ľd3�=,U#Ta�\�� ����é��ifE�+&.)��چ��@�ԙ�,
��ٖ�f���$ɺRO�փ�t�[�MJɱכ�iǈ��(-%<$Ւ�'�����f��%���^�`*�^EpEa�댟�����\���מ�F���iƍ���9�H*qTb.��`��7엮��	���?9R�k���L��ԆB�C�N�8�����uűQ��ڱwR��]�a\���d��&#kU���j1��A����4���+iy�*�u���Ѳ1��y��{aO*��y9�O�">:��WM��H�r4Y�sH�ɷNY1ʹ����n\�9�#��(GP�V�|&��Ћ���S���N�f����ۡR����z��VJ"9ﯫ5��'��k��^Ӓ�+�)���;�k�9���y+�r�8}�m(�O�O|1�����u��WQ���*�0ګud\��$
��zu�fq�j.;�a���� 0��U2B����jP긑,��,f�gi����
U%R�
��@�k2+�(��`x��GX���	�T�%�����3�Ӓ#:������B��HZ�|I��l�▓B��|B��"9M����W=L���P/���?�}&���(��Y���Z�K,�t7gl�n��#ϖ�Z�0Q�g�{�l}V:��њ��Bo���W՘�S�(���
��)�m7�>�)\uW�.ې!KтgF%w�����tb����*f{��"�"�L7���H(�w��#�Ø���IЩ"^��)�0	�/�J��e4]B �Wc�z�������'��H�S�0"̴�X�/=�.TN�=�t�٠#4#�%�{_<��o����8�?��h���l���Al����⇾��#v$=�`��� ��~��ӈ׼��?����G?�E=�����]���5'{����_�S��c�E ��K��t?�C$��蓵C�H�	 ���pBp���'̻�,���� ���1�m��!24    IDAT���3�ʪ��$���f��P9QJ'���|������USA����֦j���+d��m8�o~5�TʌC����F7���_�i^�v&�&
pT�0m����滖&Y��,�?�`������q�7ę뮏��Ɉ����: g�mL\l���[^��bg�d|�3�[��f��/yG��o�7�NoT�)�uI7գ�@ �>ᓰ���h��C�a�3��f��nl���xO��/����O��?�	{d���4e����� $+�mE�����_�o��q��?��w|���m��t)B�U|6$
2�BUJL4�܁�C�<�6{#��B⢄u��K2�n�,�3:�D��ҭI�<V2#�-��N�nj�D�¦K�+��Yh��6A�%�H·��@��|d�͜�j�1�4���C! ����b9��������������d+C�?WK2ip�%����K����21�0�@�C�6�ًm�D�ӳ���`-0%:"�J���#��9g���mc������"+/���(����;V9W�z�jp�'n�F�bb�qIJ K|5����ل����v�Mr�R�"��j�g�>B��V���2-Q��$%Wy���}j*[y��ϖ=��w���#�Q�*yV��F�~��L5������7�귬��ӱ�q�M(D��eY�����J��v�"��6"�r���
�u	۶���4e�&�� �"ͪ���{�{����ړZ�o�qW.���D�֪�x�+� �X�<+��NU����-"3�ȊZ��%Q���j^���ص��I\K��T�*Y�V	��s$L�l��)��Z,������5fE�>�~���������*���S���L���Lk�[����`��"�s��yp��Ȇ�l��<��դR+gէ�G.�e�&���'k�.�'��� _*%伌�)���ܵVj=�%���*P�òKX���sȺ���m����֚������%ߵ"��+1+�Gb,�Uӎ��*�U���\<��J%_�DDD�F3�S(��������� �ir�CV�+�˟*2�K�'�STM�L���+���=��g�/1���7���1 �t�΢'t*�Z�ƃ@�;��L��Au?�6�It�c�����A�5cN��(�d��>�D+ v�m�3�0La� w^��"�g+�F�my�مx�#���iL_���o����n��9�"hב����0�˃��^L�{���%���q�v/�}T�)-%�h�:����}0^|�k�w]��cW��9�w������ཱ�;ם��s~���k��i>���������d��2F˳L8d����ga1oQJ�Z�C��6�ڊ��2���@ffR �2��@���A>؜<�;���R�b�*�tsv�2���~��m�r�����(}���䧭	K���&�Q�[�%~�Ms852��A����s��I'x2�E���il�%���sO|���ҥ��G����k�D�<��$���d)+��qPLg�xío�������'?9��O�!��E�<��o�_yޫbΊ�$��m��� �j"Gq`�z'�꾂Bg�H柺WHPI��M�k�6P�i3��^5��{��?����G���(�ko>�"��C)U�L�,si��|�;���'��e��x��?����u�X,0�4���U�/F%�t��Z"U�&�p���| ���Z��Cs�=e<���!��(9brl;�L��Xt�d )K);�I�iN ���̖�8@�'�}��k<F�(��OƜ[kw�d/H�(��~`�e槞��)�{0��Z ���
e|�k0P�zc�J{��ӡ���v��+�(�U
���$��o��L�!�tdAE�&Yq'%)eB������$z��,c9L�P�䞦�ɱ	GX�&��uf�h�o��I�W�L���5��>��n24���cY�A�I&F����Gl�C���h��T��K�t�3}"�h=�`��I�J��zF�V4�g�ݖXR�A62?e7Y-\�<��������7J�3F�3U�X��)��gH� &��6�SJ�gG�L�ʩQ˞Z�����YQ�q�g.
t���;Mߗ{.�9/%���	�V�bݒz�k�+eNbD?/?��1�[%�Z��˙��s^�Z�?W��cۣ�D�;[*Њ���1 +:ڳ>=~H�M@�~ƚ�'�𞲃p1�S� �RJ�xo��ɱ	�]�զCZ�q�H�Hn	�N��ٌS���}�c+�߸��&h{@Y	��I3iN�3q%7�T�m�\y�9J��oT�&A��ž�D�EzMט�thk��K!���T��E+�&I�ʛCmJ���!�T�+�/�c�5j$ �ZK�`�1�$8#A팱����]Hg�Zh�Ø�:_��[ ���R�x�Q�u,8�+v�s�dA9�2j{��2ʱ9���-֝�������Soq,��:S��UUDk��)wU�����ڤ�#\c�\b	�F��GG̊VY}�c�i�  ��.d���y���}8�{�l!�=D�f���&C�e��5�8�KdH��d�\��|x�
����b.K�F����fH�Z��SK�,�$�K��1LY���9��}Iy1�_��g�c��5�G-0����|śX1����"l�F��YV��\�G�.�v�M�<_�����'v��c��U�В5���ܧ.�{�3������2���@vۇ�{MS�s�|,��G^3�����+���ǲ�L�v��w{o�����1�����7`�58���l�R��h�͕f:�q&��k��hЉ�D��~9id ˄������zփ1ϫ��贯����gG/��#�Ld��]9+Yi��{'G5�p@;
�e�?%�j��/�gU�*��5����;Q(�����^�)\B�I��������Kq�҅�|�"]��|z���8{��q��ч��g�]�>62iXo����+_�����n�o��o�g|��(�3t�����1~����I��d��� Q�G�\�n��^C����\x��
6%��S��*���^��O��q�I|��?)�����cu]<�ڭ�)�7S�ZeO��45��t���u|��O��n�#���;����n�b[�X���z�*�(�e��@�sj�I.9���N��4��  {�'��2<��b�p�~\�x['����6+��ΊA.p���< R#�ٳe����:��w,'s�,b��xD���h̞R�}�R$�kIy�VrHw71\wٳ����p��@Lr6n<�'�ڡ73]�1E^4�[\�tȕ���d�g�ɧn�$�2nH��d7�9F��]�E&��o�g桟�Q�-�H�{(3�=^޳�0�e���>�L�2ɑ!���Z�s���Q���8��dW�\+���3��@K�v4y-`>Aa�<�}G���>�I
^��u��e�(
�$L,�:T�ʵX�����H8��2E"�1��Se(e��d�������D�̚�T�G��a��wR>p�ٰ�����p(�Q�)��*]V哯�,��^+b����z�I�1�iV�t�j�G��q�c&LE���뵰��CV�h��+��vN/^{�[-pJ
��1Y��K��Y'ռ�Z�0eU���u�T���	��\�J{��;)�%���:��I;@��q?�4�7�_��<CHf�-e��E������Jm9Ͱ2?���e6��,JB�H��.�>)��ԙ�～�<M�L�������NPB��J=�����SS%��1PǷX�B(+(Vx�3�� 3I�K�����	������?HS�ha���"�}�ٷ�qQ���y�|����@��V��{�1[���A��J�lU7��W�M���%PvE4շe�P���=�=LB�G�>7ϸ����wTg!�6�}Ɗ�hQn���֧JN��9)ޓ��}�=�U\*��48e^��i�����(��K?�?I��p� ��al�V5!��8:߿��p��V��^�z=�����=�/NQ=U�����Q?:��bd�pH#�R��e�U�m���g"& �᳡�� �j4Gk
�S.���1u���M��I����2v�R<WW�Y�E�)��p�nL`zәA��*W�����_��qi�]�)s�e,S:�v73:,�g{��É�0&�!���
2Z8�c:��|3��p;z��fê�ߍ��^|꾻���q�u��_�����ttWK��M7��؝������=���"�����Lb�����V˘ϧ��k�N�t�����00��u��-�U� `�/e%�)xHd0��2x�F�`d9�3��^G�/y��ӟ��r^�z�	B���H�~�{X�O/����:0i�ͫ���2Yn~Q��0�Ty��Ϟ��r:�Qt�Z�%Z�Q��96�bNm�l:����a����t��fN�q��8u�i��;q*��3TE��
UI^R8g��d�8�����m��W�:>vם�?���o�:�Ri�3�D<�^����ǲ{26�I��[�s�)L����E���q����me)�N��"xp��f��}�蛍Ɛĩ�Q<��k�n�����=:n��Gƙ�o� Z��<T�q��&>9�_؍�?�p|�OŇ�/>ya?�ݘmF��wي�
�^!�>��L�L�����a��và�#�S��%P2$'O'Td&���; �Ǯ:��(���/CIx=Q����@Ίke�t���X%�c	�g�e�)%��RuR��վ�P�U�f-I8��� ~q@$��
	�C<�A�cgX�%0��w+el�Q���\�0.`B��	%z��'���c������x&�e׌|�ן�5��ʄ!�ʣl�e]�+���V�*��%��'��F�ژ�iU���?�������:2#�kqh=������;K۔:a����D'+Jr��r,�	���ϲ�W(�q��=:j\T�e���;�*���9T����{�Tko��\YGT.��Y�sb!�Q�ld���rE9nG��%5s�5׮�CL��3{�����^\�6wr[U:z[%@����L��G2�aO(�5�(p��z��ïC�_S�[��@�g����-��n^Z���id���W��2�0�d^�T_���S�X�~#ټ~}6GѪR)����.��+;0�y�i�:8Ϥ0;���sh����t=�W��3Q��ɓz��W�]�w�T{��
�DD���ϴ�Yz�����9N��Q�`�Τ�Ѵ3�ⵖ~�<�H�"���b��^�y�Ö֮�����-dD�V?�w�!O���1���N"�N���mp�!�G�fd��^Y�Y�<�R����o��2�-k;����^��U����9G]�J
=�$)�����q�����V�r�'�����G��@<8�y�]�7TM���&}��_-8"��L���mMb=�ǢEv�x�J	)k����QG�^�c��r�( dͨ�P"�%����Dcd��U.��y�m"��\(TLg����̯��z#�7� CB`
ٰG�p�Fs4:�2w� ���5�r��a��h~��?�=;`
����G�W_��ٲG���Q�����%���m池�%�.��^�	v��6�x��gm�Bu�Oi.�Y�n'Ƙ[������}*>�;��_�����?"x�du�#�(���o��8�Տ�`�S�2���(�@�ɜ�t6;���~��l6���4�Ȓ1�u�8IF�o?F�IC�� ���!NVI	w&��B* ���◳aF�����8VB�mmO����Q9�-����0�ft-U�uay3��Y~�(�W�tS����R>]��v�\;�����	ʘ�2IS8�9+�l���K��<�4nh�;�X��S��.P��9~*�:s:N�>�N����vt���= f��pZ��Ø�KV�~��x��������b�����-��� L���/�Ɵ���Oc�=������� `*��p9Hͦ����7C���/K%�C�$�����y[�M\sj;�=��N������������f��7���cwk}�U/����1E���* "��e gv��)�k�)AP:Z��ve����h$ ��CS������t)�9 S� �p�ݹ�d�ǃXlV�4�d�Q�B�Ny�U'��5{0�{d1� 3j����u2���$�=�x(Rp�2ऋ��g�|Y����:zp��!`/c3_��pJӉ@)A-܈' �ʘ�$v(OS2�D Y���3�g����F@5�m�F�^�J&�"�D��	���@�
�@����.�X'���{�
��"��-Qr��_�K�����TM� E��)����$vm�i��Lb�1�`]�\��i �)�2��.����LI{V`���(8��e����q/�U�����_�ܙ�ˊ�\']��4��Ƽ>��$�
�U�iJ�Hr�5k.�24Q�M)���La����E8�1��ʙ�$gy�2n�Wz�ve���F������￉S�1�&�m*"�v�^����+#W�٪Jm'R'�Z���ה7{�+��dN7G7Xj���@��+�j�pũ�SypWT�����cI�]Em�|��Cyu�W�Ǆ�Hϵ�MqY6�d���g�DD\ه*�ї������2�i@2�H�M���L5�iWG���vO���SgY�u��Q��vQ!lLb�� ��#��DITq���� � q�|���/�gCn��R���b��,�f\JW]�0��Lf����ĝ��� f��E��6�������lӤ#�G�~R��"�� d�X�1]��_���u���m��i���/�
��k���-���2Z�#u_�;��H�
H�tM�Z�0�� ����̬΃��$�(��vk1&8չ��:�j�D2K�tb���	\u$ų}���I^���0rD��߆��9	��<L���#)���� �hWZH��Q5�%�SGb9KΙ�B�=����ܴ���P%��0�E_Gw�*����F�+?�}q�i���+昶�?|���W~�����R�L�)��b9WҊ~��~l�o|c� �p�C)�=��Zu�(�!J�mֱ5���`/��c1��T<���O�c?��)��b�y����X\홸��Uq�铱W*Ved��@)fa�r�,G��'��a��^	j�W��:�9�k�P���?,gV2�J��2-�\��n��x�SP/",��FHg��><ڤ�=H�@�����Ĉ9���E�J���JP�kIyX���`�U[U���I0'
I��lD�ɾ(�w�6p�Âן�ff��|R�\�]ΨEE{<�D0��} �$?S��S�dg�hC�q�?��>~o��e�-���^����O����&���*h,$���_��x����R��oEw8�5�� ��� �y��0��Q������~�Ys�'�:�X�笠vV5�#|Bƾ�E����K� 9B���!��b��� �@�1� 2�f��j�s9�Čr_!�ˊ+���!*��ˆ�a3�*PI�`$� 0���k1��N��Dt(Y�|�wI|c���X��{����C=�="X��%x�*,ggj�����q��H	L������`�]����=m�~0� �[x�1-�Z$B����^�g*Ҵ<�3Y)C�]6m��-��k0�S"#F_{O1ȣ���1N1�FO�$yL�᜘3�Q�:�fj�J$ܳ��=�Y3�ѥ6s^��
�\%i?�e�
W�=����fIB�B*�H�	 �`vE���+,��1�-"v˭�I�q%%3f�YS����)g2Ѣ���Q�[#���]%<���yR2��O"Pyq�6����յ�Ur'�u4����U4v�d_kş�Dk��+k9�μ>�:U�d������U:���gR�Ů�r\���hݬ�p[�"N~}�Ԓ�u������$ �7КL�����\<�i�}m�ڸ���S�ay���җ��T��:�A@�q!n�Xg��k*QψauW�@�n@x/��V�s
�6�W�ȳ,� [��篶�B\��\<I��Yk�xſ��w��e��C�Z�ʠիi +��I	�$<#�x��x�l�ȯHJ��鬋5M1��    IDATg��Q͗L @��3c�L�d���d�m&�er�C�Ϣ	���t����nR>�_��_*����dN��`Q�y��jS����@{I#i����j�&|�ܔ�p�>D�(��	�H��|x=��JӯP�-{��=���B�|�a��E!Y���Lgg�v�|�0��.rd��w�=�Nc���pN�H�o#�/����G'��.g����1v)��|X]7����g�Qș�cv���P�@²���%�<��"7!�*ͥM��úѨТm	��`���!�)!�A�)�.�L�H���̽_�VEz@ʤ*��w���E�W��>��b��f`�q1��w�/��5�c:[�]T ��� � �����L3K��F��:����~��S���x��;cz�\<��S����L<�;��L�N,��x׻���G��ӱ�5��O�ӧN�d8�c)p
6Z�|"�Ұyo��QW���9�, �����d�X�R�i|�or��}������Y
�ֻ}�W�F��G�/�����*�V�,-�������u��ۢ'߶�+_6�U��P��֋o�uf��^JK��H�H&�_/%�|�¨�2�õe=���`��ɤ�I:�5:q���q�m�����O_k<|�R�/��{L����x|�W}i�ѿL+�����?��~�[c=��U��pB+����avD'D�M���g�	�Nt�]mϊV�wKK�>�,��L�e�o��$i��HU~Wu9d�U0ux���V��=r� f�R"��x(�&�10�cЋ��VtG#Z�����$P����[��1��ǞVL��܉���)���9S�˹�Y��0�k����!���|[��>RTmi�Ι�c_�d�q-��J{�tP�Ve��8TK�љ-#h�4O�.L��uU!��N�p!Τ��7�
��%�*���!g&�I}�{��_!�o��#�H�3-EWz�*Å���?'��٥�(� 268qg��3�\	kf1�e�}��(ؐ��.%�NHR)�{
��f�F�N��M�Q�c����|
��K&�T�d�7��e�Rr��d��Y��UT�4�AsvEȰ������Ӫ��}�_lu��#��v��X*}%ح���g�J���u�:�{
R�QT���Y� ,y��^��pe�G���D������Ȩ��I���j��kK��џ�O�z���*�P�d�<���M�&����:A���]Ngw�	v�R�a|5���Y�*�@]r6�2p)F��v� �
�
q1�bʗ�*?�\�H�s-�:�|+�Ic�$)Db��`�=�g���:+S24��	�x�uν\)+�dl�^+��U����nwL	N��#�=�b�r\�\ʹ�
,�|)��;LyƠ'0���J�#0���Ead�jU�c,͵�r�@	,����f�Q�K�v������ۄ�� }�zV�lgF��e"3�S��j�,oE�\��go��G�i�rk��k>IW�B��S��J�3�ەG���ʬ=%�3�VS��?�Sh����>���26�3�e"G@�@Y��W�V�rT�i������$��]{Q� 9�y��S`����x��R��y�k�M8nf�X�?4�#��D �Ui)��H�;�:�9����`�ן��	*0�@�y��;�
כ��KiR�*J�x�E�L{���/��G����M[`�'�7��yu�c��U��-���ZSj)f+�+tR���$�<�9H�����X��� ���X�>7?�������x�ՃPZ�
�:n{�����W]}u�r���d;�q\u|'����U�5� A=2FʊU��H	���(V�i���g�P�/�K�j-��NPr�*�5�ё�X��g�C��˿�%�$Z+�����J�>�˛�̍a`T��S��g�=+Y��S�����+_#�����`��}�Ya��@-h֟)�e�k��:>�����7�-�������#:w�����0��ω����˿8�=l�^L7?���:^��D���vP��d3���ل�U�ػ�ɉc���*d���J 0�ɗL��I@Iz!�l��2^��4#{�\� 0E�4H��ېu�"-�+���\L�rfN�?�Z�Ǵ����k��x\��������!pC&2��G$6��u����ؑ䖽+ɍ���`�;]EV省:���%��Gd1=���ؐ �?�z�YQ�t����>*�8t:�et���D*���tU��X�o�[<�WJ`����hrVi��9��س"�U~8oe�uO��du����a���?�-Sjü�{0����kHYl�����N�����=�$�ɗ�5�E&�����Co�|����{�Gs�e/%�`����Ĉ�}�����N��֊�N��h�z��3!J��ϖU���9�rC�<M6H>j��<)��+y	�s��p��a�W�L��
�T���aW2�- ����z���se��= T"	@�O3Ac�'�G��e��t�-��ٟ��O�[ME��d)�����V��u]��;g>V *��D���S&�	����e�M�]�N���(��Q��V�DVd�^Wi�%ܜ�aV���
;Nn����=�9��T*�x�B��I�zU&�,��oi��ky��	�ւK.������]�W����ܺP��P��=�£�^��O7�:���Ƴ�Zq$�Ds�����R�j�����[1A�T72X"p�ʸ&*Ԋ�� Z���$����.�p}O�{_.[�H�����/J��z +�>��?[�A��R$�����i�>o�?g��D��-�g�x҃o�����+)��[��o�uš������+��:s��
+s*�
k�i|�	�'6�r@bEd������W�U Pi��<d��%L���7��Hu�\��ıo�th���E�y��v�JfE�:v��	9�e)�u/%���.��������'aU*�̃D81��A�z���P#��p7{N�����p�A�Ԡ+�ŲbJ����; �DN�����.�?;�����k*���z�,TL_s۽�/|����nl �p�H萊�;��ioN��@Iz���0#�:��ѡST}����a��X잋��x2^��g�A�G�o�w������a\�|10���{1�kO__��_�z�E~���������L؜�<7 7�K�:M�@KP��1ٻ|�
�ZF���j2�M%�RY%E�]Q���*�F�Ӳ�N.��Rill��{��r���ў���!�]��a�d�>C���ת�g&A�յ���|.��<�q��n�w߹�Ї��q��?���.^��b�a/��x�>7~���C|ѓ�=D��(�~�O�/s��,{2L�"���h���e��ՕS$�%[�ح��JP�ȡԖ-�#@�����i��\R,T�C��j��t�6��q7��|N�,{��(�=Z��:�d������yZCTL{id�S��Y� ��M�Ә]ڍ��!eQ�t��U1>���p�E�M3|H!�;���*���{��"ub�5��& <=�l�cEo<*N�g߲:Y�^E}34鯣9//�|K����@֍�^`咨�
�����`]Z�H��~���	4�L|Pؤ@KKU�ϴ�Ҹ"�������*Fa�VeMJ�Dd�sS]��à����f*m�!��5�K��g���I�i��ѣ����[�'��Y���~��������
(��}$s��������G��C����z�����)�0eH��'��$ݬ��̕Z̟Il�
&�YAdRY�̎�N�D,%��
��I��S�j�9���3}�.��T�}	}��&F�VB|~��mV�̴�C���|gݿ����B��n�c�g���um�a�d��O��c�eݐ�g;O����7��1��^H�=� W�
�%�B��g˰��qDh� Hi����75�g�s��j�?d݁V���h��cR�@�5�yo�>��L3.�O��W*7��>����7tV?
d�w�Ʌ��7Z��*��X��+��v�����$�T��	nT����1���
���(s�1�g�v�Qn!����8�6�V��x�8^���7��Qm};���@ғ�QG󣀺��0��(����*2ᣊ:�z�9')+����L�?:��rp�,Y�/gE���M�=����u�Z1�f����e���1�J��qLY��r�����2l��6�b��߽9���m#=+��z
`ׁ7�d�q��T�^cK�2�*��U�b�C1O�E �0C�1*��~� \��8��#����L±��y��Bސ,/�s��b}�^o�=����j7�;<j�~l���c��b�������F�K0?:;"�S	��NL_��{�����r+�~�2ّ~#��_�S����4�QƅHnoU��$��4M ��v��x������=qӣN���W�4�xQi)G |S6�;����e�����c����D�'?j����2�f�#e5��C�^L� t�\4�}mdt����ff3qq"��<+�鬒w	�G������J���W<H� �R$���ǉ����+!1����Im��
d)q(�i�A��d���dᨯV�&¦_T/�0V��)�K�.�����:��U�;w!��\<p���|y7Y1�LF1����/��{�W����p�u"~��������l]�5t�C�V�P��`["����b4<��3�s2r�g?��(>!��z�Xff�*%�]�+5�@��S^'�	�YM�$�LJ��%6�ϛ,:*:�Hs#$���c���5�9:� q%��$#�M,c~y�fB��N��gN��bPy��ROx��,V1�4y����cvy�f Fǎӄh2J�P��=�r���18���XB���#�6zM�\
0B�d؏��m+�>��g�G�ھAƾ�R��*�;�n�A�=HiJ�}��nb9�2�v�;ٷ4N.�v�	{�i�/�2��ՃJ~T`��_jI����]�r�	�R�H�.����IF9��y?�>3$^i�b֞	�{d��3�����2W (��ɞS��gA�ਭ�	��FV` <������bgF���a���n휓W+\�	0���-���+��
E�f�$�87����E�\��K|VB��c���=w<��m�9G=�=U��D� J��|<yJJ���!�ϟ1Y³��[\1J�,0R���k���8�oA�����7�5�������7�D&$s2H)�(Z�V���ZZ8t����eU��XmW�N�(M�8�ZN��"*8����*�If���������Xk�uι"V'������7���^k��v9/<�	|���*O�$�}�r�v�CfG�+o�a�w���8.Uc}�}��n�֨�U0��BR43K9bD������BzZQ���$eu��Q�u;k��AW-K|��T� �ҲN�kTP��j�����e<���#{����W�ر^**,�_��-�<ʞ\0��l��B)_�D�99��V~V��P"^܇�;�3�sĝ�t�1vZ��Ĳ+�:��/<o��6�Е�2 ��}^
�G�+v�}ڴ)�B�~�Df�cM�
��|�~��=&����N�Rߠ�+�򾣳����(�R�$cYө�, (���r�����c7��I�l�n��<����.���T����8�� {e�⟕�B2�Ц�Ơ8�8���>9���2z+��ce�4��*$��h�<u����YE�K#� ��Ȯ��� �=�S�z��Η���)��)0s5��M�����)
haj�N'A�8�D'�c?m,Q���"0��v�g���-�������L�ؔ���M�n�1X\��?j/����'�6�p�t�C�=���~�}��/�ոW�-���ڙ�}_PE�ᙬ"Cw�x�rd�<E &o>���k�����]%0}o<�	������mG��6J��2p8�q�V�D�<6����Mn���!�~.*�V��Dɻ�[�S-���*�Ҕ���?���3��?='*�TM�fr�p
f9��]mӏ�}��nþ����Yt��l���G{_U:䄎�>���]z���=�C���x���}����C����	���u�n�0��夗n�}VN9�4?6�p�~�K_K`�;� �pg0�#e�.�aL
�l�%��p�@]�<����|��yn��_�%��� ��a��<R&O%!ϕ���&]����v�Uq�֏���^.�ۍ%"�h��	ٹzX1��_�有���af��_��ق�Mz�a�q%�Gj؇)* N�%QF�.F`g�8{�j,O�1����;< P��!Ը�W�8�Z'���M�EV� [��^�5d�
�<�ph��c4�}���P��W�I����%l[�;|W'v+���=�1���6�4a�YH�#3���'Iz��w���#"��Ε�WI�~�ߓ�Y�HWO�����F�T>���6������x�M1�W��E��Қ��O�S�gEI���m��Z,+Z	.�ge�LD,��(��R�T��L���ń�y%�� !t�RN|䈂���T{4��˟�>W'Ym"Yj���P�?�������$>8p>�Ɔ\P����yXQј��<ks������3�>'�YQյ�*���iRb\J��0�e<M)Y=�j3s1~�X��e�5��z���TX5Ӝs�^��uI9#,��#�d�����)ȳ�~{r�X��޹����3�/	�$��q':���X?��#�Z�t���V�@W� >٤L���)g~yNR�(�j��x�6UԌ���˄O/maj�R@�N�P�D���ɴ� �\�do�ܛ�=��+bN>IN�����n1a��^��晾.�U���!I����x��fEE]�-���T#1ο��cߩ�q��ՊS�6kΉb<W��"���T��
�Y�4�b����B�T�Se�O���l�)�ᝁ��f�Z��� �^K2��C��"�n�ۘ��Cn�֪���a~�D�gSW��m�z_@y�\�E:�Ay]H�E���-�+ ���X���8_��Z��O����'8�˳�E �z}UM��OTD@ҵ<�XA/�6������Qy�X�i{y� C�;�u�r�r�X��$Q����q�.�1��b��O{�(�˷|y<��0� ӗ�Z��r�D&��m@5J�1���):m���� ���r��+�gU���m����>ή�?���[��~���<�BL�J�
:���{W���E���X-��޷�-P�|����#�JV�Ь�7Xna 55i���a`2��=Fq?����yq��`=͜?P:	Q�u�g����{&�_�
�]a}�>ekz����ר���j�t�ǒ�g��(ϱ�%���:�r/��԰���W�x�8Q��Y�a�|��h-L�&����ї�.��nt+�[8K��=�u����Rn� ݰ�5ث'�RGKquU���sB��Y���}KɎ���=�y����ٞ��rqֵ�X	\+e���V�N��������IHM@@�`ʃf˞���������]�,��O�Q��\Qā�.�+�y,�^���AsSG�;:���"�gC&O����)׆�3R���($����<����<��(����A��n���:I�ﵘg(>"����]:�	���O���}��,�I�|ޅD����ʌ~������Zw��Ye_<��q�Z
�
y��HА�4�߽5^��	>��TA���΅%�TL�[+�i�騙���Xz:SJ�� �s�&�Izk �+���]�-�N3W�Ě�`�m���F��1A�$��--EI�a�b;�6����]*,�}��+0m��(UB3�SWr��m�̘��夳 �*!.�1G��ߵ�*��yi��|����Z[����ė��k���MS�y��)!+�ձO�Z/T%��ʊ��@6�	d��Z���S���
)�kO~ν\���jif\�4�rEB�R�+g�+b&	�D�� �/�>�Ϊ"�@����2W�M0�f�un5�1�j�r�9��9˺{j�T�����Kb�V"\GfT�IfCt�O�,{�?hL��_�8a`�X�1^{���1�p�{�*n}�x    IDAT�P�5暌HB�ϡЎ*���>"µ����1�2K����4�a�pt���1���J�G�$�%��-"3j�� ����6�\�i�p�ٖS�yͻ��`��J�
0G���Ŭ�{��SN�`��syq�G�4[�R9���!0x���c6�rho[mbUI�k�yP5T; �6��nK�v��x�]��7�!8�)��)�&���b�e�����Zw�i(����w�v(�
@ֱW(�0�%1#�f��/$�0E辶h�*�{��F#�;�*CTf�0�Liz���~��E������p�4����)F��|_VF��D���m�\�� sLp��}�W�=�b���e��o�@��e����Q�6()��H�T ���Ka�������U5��)��;�ɩb+��f���f~5:���^�o�?��▣n��X�����)�/����v��I��o�&.]�O}�3�ʭ���E�>� ��4!��:�\�E�U�6U[�v�4,\#�Ց!f��?�*�Q�]9�>0��-�\?����#�֟_�Lj�C]o%�ٿ`�k=&3Mj$��O���l��o�}���DY���β"}n[s�'�@��0dY��?���t�/��������o��r��HC���+�ަ$�$X%�,s��;�k��E��җ�3f��Ȟ+&�!�{�c>,=��6��
,�@/	s��p��_���h`�bpt��i�+��`�yp���@ =�����b��������� �恐�ayg�/E�{��-�x�݌�l��Ð�/\�ᅃ�,;����I�SIљ� �bA!�S
�`o�K����{�ؠ"���w��ՎgA�c�3A<*� �8�Џ��vbu�P�ì�����8�y�k)hF�@�#	-d�\|�*��K&�<�"��c�8��BeDk�0	����[N�]�LR�������}Gӗ)�V呞�?�P�O&Xɪ��	��fQִ�)Q�*��<l�ȉ�pXu5��<�x�	�-�W�[��|9VF41U�4c����Ug���_���VE��UMj�UIg�_���2�ǚ0�=w&���R�J^���kȄ���Ȉb+�$�؞�0��>z�:��|�N��<˾��cS�H������ y�C�9�̥<���3-FBC���<�-qV~���z�Y�>'\1U�^ﭐ5�J9�D�w﹖�����nS��Ds�6%��Ǔ�#]R��:Sm�uj"%�4����=��O��qC�F���e}I� �?~_抜}Z�v��l��gV�["NkOk�.��ۮ����RH��ɶ�/�����D)骻۵�;�0v!�F��s�  �m�Y���
0�~Ί߹"��0�;�Vb����@�8�D%�C�j�>�4��#�2�օ�2�R�Hz����r�$�l:��^IK��K�7�<���M�8*�,7߱b�����IXkt��Đb6�٨�bo�L�D� �r��z/a����'��$KkM�tW��Ue� ��:V��~6��bż��YEw��>�W0wD1.'�p��:p�l�L�c��y�gI�JN� �N?�P���-���J7ݵ�tE�h^*Tdh�����}��(=�ivF` ���X2�q�)�V�#�3�`Me�Q�蠨�i2�������Ϣ7W����ɷ��q1�:�z��.��ËA�Q��A��e/^
��
��=��%-{�C��hy�fe��2i����4V��qr�q�mG��gd|�Ӟw�qKL�j����>���z�Q �Y�٭W1�q-���o��j���q��<'�z̝1�܏,y&+� j؟���
��'j�(8��$���o�J>:JE �aӎ��4���?��d�`��A�1�F[�*� ￲�����kn��^lr��RC���6��Ϣf5M��������Z�5�a�#�ߘ��7Y�;:8�.�dv��j�9��c����6, @��:�=D|���L�������b:[�h|@���՚�*��1)Ÿ���s�����b\�G���%"�!�ǰXB}�XL�Sd*�	K���Z�ؔt;���0UϚ���Y<8�ht��]VLL!���}�)�$0E���c���CWcv��~|�=����`(�ә���c� ә̏�3V Q�\F�SSH���¶S�Ѹ��䮷�'�T� �p.�XK �+����tI��W����Ѧ�|�~:�uV�Xc�X�쐴��[b���yu�g)C�r��f3BV�;��Uݘ��+�3�[��IN~-��2�sΠ�j��L�*���ѕ��l�&ʮV�/)�}���ik�&['պ���	z)�.���XO�h���9�|C-W8���(W1���FT�>y�z���	2�)H���a�ZSo{L��7�&S��=̱J�Kf(�.rR��������{U�i���zS#u~z�#\I^�1\%���":�6:��;m�8�f�T��d��=����ڄ�S4�\O���N�\�c��܄����3�KL�%xd��^:�k��f9k���U�'��M Zj�j�J�����n ���ẶoEa�:�IՏ<?�:Mfl���/L��BE�� G$De��+�)���Zn\)��R~g۩h�{���'-�"�
Z=��1c�Ⓘϫ���F�}bO�$ R۾;�����.<�4�=��h��zkј��C���J������Uh\��I���q����B!���9��9����sY�=�u�佊)�����=�i�E�%�pt(��C@^/LAp�*;bG�h*ǫ$��$(���sh��P����ť�ddB	��� �Rܪ�'S�"��禍-/�aH���&bsz��7c�ZG���E�����>��[���q2c� �Q��!%��� ���2Zc)Z��l�ڮWeVTl��y���s����@�������	��rE)/d�p�*�����BB�=� Lq�A)�����0���Y1��7 ~�富� [+�����]���:�c��N���9ύ؝�gZ�B��v����flWS������.����x4�\�Lim̹B6��?��0���)����$&�q<�'�3���x�O{��ʕKqt|�I���^�b����%�̢Y&ANJ��K��2��k�~�MS��jF���ɇ$���U��!K����x�n�CN������9^Ԋw������g5,R�^�F�gY��I�����,Q�gɣn�"8U���,lm�4+Z`��jg�Y|���{��}���N�b8�w���r%&���L&$2ƣQ��mW3�Y���#)P/Vۈ��<��x��Y�����������0�˱�tb�5�(GZ(8������pq3�{���iJ�JV���]wv�+�a.$�Q���ȣ&�T��-&\ihr>EW�R�UIb�ۊ��Ã���Nll ӣCI�{ꑀ��$z"�L��L���k1?�r�B�[�iOfB�SQ���(�1XnY1E�G�*bR<��˗��1��A�-�ַ��4��&�s.,�1�fGKIm3�C�#��1���70�5�ka�D�<����1!809�,��.1�F�g �1bK�S>%���3)VNl�K�k8g/���"�"�n��p�U�>N:���ln���\�e�ɳ��4߰�I>��Dە���$���+/�$�����HtJ���������O 3�.��@� �M�
�dCw*��ڊ ݪ-�H���%+h����Z�Q�5~�*q�HeE|���
��Fw��3��'T̈����&4�m{�\YI"@ϻL��U�@m+-\N��	��\R�1���A��%�n�IК�rτ%A��-T����d��'��t���z��>S�qm|�w��L�O��,"n!�DBZ���MŪ���Oh�_�5IO�	���Q�]=�5�he�������`L �J������(4��D��\3[=4�f#��X�*�j߿����5�{ȵ�p��?o��BC��s>�6���虜�����B^ݣ��j����橍��K����gG��@���e�R�
�=�9���V��Go|\����r����>[��A�˯�%���E�r�|V�\�s��=����]�0�6��4�S&��lE{�S�-IwҎY1� ,�pJ�����0)@��i��
�2�!~�u�=�D�dU�
�&&ud�%����3�b�)f��rz2�/�&�b��4����/̉� �P�����
�4q�^N��I �Z@܅�3Ti�9G�`��
2\�T($�I�����"�z�d����`�Ċ)�fW����Q�I�H�=�R^��h\K��w�^j\�\�b~䟮�
��b
)���U��]?vp��HZ��I����T%��������!�ņ#�D��|,�j��w+�+A��r�%�e�V��*�C�O��&�.����0A���1��f5�9,�7�{q|4�+��c<�ǣ�-n������G�c{w\�|9�X�]9�)`��I��6�AV���K�w�'�\H�B%�J�͢�%v;1
D�F�888��xR�>̨a1�,0�h�e�p4��st-~�}�|0X��U,���"��Ә����r��)\RW���Hx�ԧ�Y�K����[�y[2�@�<���3	��Z�1��H����]�nH����̮�-T�V�A)��VJ,16[�L��=^6.h�5N����g��gH9����|�c�� ֽ���hzD-����~N2�//�/�~�� ��:�Q��~V�ә��܇��J��aΖ���Y5��!Oi�P�X^�������s���e߈�B���(��ȋ���Gt������Rʋo@�<��"+�[���!/>Ha����b�ڱ��I7Ê�h��l����@��!+�f
�-M�0R�O�����Ѥ��`�G�H߀��u�=�$�}����*�������Y�|M��������>N{J�"�yDd`�c_b}`?��V�W��1[�T_�բ��3)��>�kufo�iϲr�X'���I̹�MT��<��qo�{e�=g�n��k�&�y%�T'U%z����:Wsa��R z���� �����N�c��C�/��Me�Գ�Y�J@�@�=���;?_�,��,+eoM����O=$WLO��t��!R�֓��2~5}�&����t�ڊ��y&�4sXd%:X��F~J��T����N-����uQ=-𓔽3�?-�����)�Z�Ǥ�W��Q�%Ξ���6���4�3�\�n*�\�ǝ���}�5�@ĭX?4�ɪU�^\u��U`��sϛ����G"N����f�{���KPK;|S��S��\�?�&])����[W����f��FM�%�-Ϭ�*�1ǋB@���|�߱�cG��0��jz�R`e����Zp>^�����
�j3Z��Zŝ޴��IiΞ@��=�`��ż�_������}�2����_�l��;z2�+1�k
�O)7��DfԽ�j�4�6�ӕX�LU/�zsSڟ��!UYj;��Qb�H��u�9�`H�@�d-�D8I�y�h#��0}ا�#�as;�Ss��_;0��3�Z�Y��<67��].	N�m�:�y����8�!T�H��C��n,�T��L�n@���z;z�s�{g؎��􌘀?�яc�9�la�w+�4yU*
	�ŒS�����/��O&�E�r���l,�R?�Kv���f�t�'�0����1]�ֻu�b)�[���+���8�̮A2�.�4�\���oĎɾ��|�D�G%Ԭ�ҝI�ً�I��

X��F�솷[!v�J4gbD��-� ���� @u���*xN��rq��I,�X���61�X��f`���SJ
����@O�O2Q
�@�j�oE,����L���Ym���p�Dόd{H��,�X��G�:��\ ���ɑ��Z��V��`�o
�y��?2a�L'�����)疤;?j�S�s��l��wŃ��,��j�I�h0N�%Ɉ����9�x�A/z���0�t�W[�aX`�
``Z�L��y�D�s����akcF�p�>���vG��d������<G&��G��A�#�iI���
 �P>'1�S�u��0��K��t>4չ�ND�k��G`�b�گضܮ׭�+��1��`U}�It�x^�<����9��n7�x�g�>t�O\/�%�[/�r
�p��c�������� ��Ѽq�k79n[����>�N[���P���2���{�4z �kUd�dR�-�:F8���r��'8�$%�s�S���|�bMPJ�c�&;�6>�E�`[UO��+L)�C��C����QV���+�i1�Z&)e�UV��,&�d�WCa��X��D)1�a�K��a���l��Z�<}(����v�����6�mz)�\*��g�֌�p��2�=�	��c��*�s��$�:xh	��2|5��,���5�~%��ؤ�%��
���Xg����G�@���S>�ֈ&{M���{�$����jYj��R�����/Am� V�0�s.��xT%�N�|�,1Ja�Q#�I���s��d��
ɵ�J˓���_ǱY��Vʯs��e=�	|r��m���|)�efuL��U��W`�%0n��}iAH�,��&�z���F�.׳π,�}�	�u�gpV��P��g�%Oӄ��#�m!o�Y�M��񢌱�E
�0���$\�<�W����),��~7(T6+���~<��J�i�[��z������k�D9�1��󤌗k�IK��c��^=��Pد�:����j��{^bQ�%��u՝�#��B?��{�:O���J�H#bgQ�:�YUK��!&��[�ULI�����0�?�,�P|M��s3U@ev�0"	�4���j7 S�g�&b���`kO'�#������x#)��Y�<`�߃���il1�y��#�Y�������x㇓�0��ԃj!�����n�_3d�T�ΦӘ�Am���c<�#�7���g$צ���bt1�E=��g�|;��b�A?{`]�ӓ��3�����\�n5��v��zL�I`�ޑ/�0�c*`:⸘MW�ot�u�7�,*��a�!����Q�ء�k�YMx�����vފ]�8x��3��c,2���%�U�<�`-� I<��(�c+����Ի56f�.�X,f����s	��E�0] �r���1��W��=5ܴyr����{�M�
���F�p����A�<�r������m��լ<��^�Y�4��=��JW�ǀg���<t�x%�ὐ���. T��H�Ja� 8�1E��
��3�mz���Y�s�ԍ�*�;%yf��B$��� T7� QR�M`
�ߏ�R��XWLxX�g��B�8� c&��/g�B��`އ���ߟ���%�|P�1��(+�\S�<�1�-M���yȥ��Q�	�^b���Ѷ����I�< ���G/�L=�Ҭ�0m�n��%#��v�cͶʆ}��".@�Х9昞|�*�Bӕ�� Ʒ\���MSʛ���;xm�N?F���S�����<���Q`J��D�^����-�L����69R@��$���Wz�Y�4wZ�8��&f�9K�p���Ҭw�C	��bX��,�c�����"�P�{Sr�꿫��'�E��R�(�d�6nI6��̣�IuI`��m����Q�W'�����
;;\���+NEj��:Nj�h&��a���i��>~��Z���,�w�g_�y�9o�3a�6����+ZJOA�&0m����0'J���:14eD+c��"��_A��{�{��ܧP��.\�l��R��=%85XV��J�'��-"�DkV�l �F�$ܿ�Oy��b�]�f�p�bj��M���,΃�	��YSq��wEQ�W��i�[+F|�^:�j�Z+R�L2�<�C+��iE&ǭC߹�}4�|��^��_��W��qU�ᦪh�Է,_�%�b(�^�ՕU�U��q[�`�Ѭ�������D��g��%�?������βgM�r��A��=�64�*�
6����jtݗ�L>+s.�{�; �R[z!M"����k�^��\�L�f\.Rf��6�\�נ�    IDATU�#"&�5g 8@ǿS��5F������~����o���^#4WG1�j�RD��W�_oR�Q�a�R��Lm3���r��:�0�1S��wX@(���>�CA���
i�ӽ�iY�er`�v������:Z�g�Î�� �K8݃yin	�
r_����y�HYo��3��WСZ�&P]�}���4Φ�X`��f��8��r�伊}ȓ8����"BDg����b���i�Ҳ+o���;������T���FR���a��?Q1��;$]��b�kqu5���T��5 ��R�E,�	�R��ZJ�D��X�ֱ]m���%֔�q9���*�E�͆�G�8pӬ.zA3y8 (��� � ���SA�$�yм{<�$�ˬ
���,�[�u0dc0�i��@VL����ߚ��}DԐ[R*�o��y|�8��^c"�h�d>�M	�m�C�?|7m黔��s�o�σ$�$�<?޻�嬢�A\�+��'D���{%�a�O`�
%���Ug2Z�W�ѧD�d{ �?��,����o�њ�.�Ұ
I �����s{�D'K�nf�3T��2	�2��N �� �ǟg��An�]HpBM������۬�&0Ux�w~n4C�
~/7omhU[���4�g`�G��J��ٖ��P H�o�qY/E�wR���K��L�R�IW9�H��&7G���2^TLL��ɻ��>2��^��$&���\�����Q��9�A�;BL�9e�)*�x���$o��wF�X��`��ļ&�,>"~,W�>���l�4'**��&�}�	A�x����8��i��F�ͳU=��ng��|���e�jK���$�j�y�0�1�$�oA��%�q��g���,��Wj�5'�I��숪��N$KB�x�1 {	�I�X�&�x���$,���I�2���N�t�us%%��Z��D� �����E	@�p�'�m�_�@��i��NIa.,�ܫ�8g_�N݉%1aRX��Mf�Ա^�AslIƽ���
�`ky�O��s_a&u+@�7���=�me�|������,{�����7��PZ��U�:�x�&����������L���i5$���oӌە(��V��&B�j��em�^A�$J�fk��-�\6�"ӡ:2��R�߲���7o؎�>�n��cL��yC1�� �9UxKΑk��B�so��.�z�t�eN9��iه��@��GY��/�u��ZO�,��)F@z�[ I�B�bA�]u�� ��d0��k0����Lo�Vly5���o��_���^P����~��?e��n�̃�����~Q�خ�J]:�l�	#�}(ش�*���R���$��+1YI;�;XVS�Wzf��!��U�F��H�R�d�;+��[Я�»�8c5�&R!�Z��������t2�*��n,�"�A�rL����`���`�;�ԁ�UlN�����(�5��f��O�#��%āh��p��)L�P��GcV�Ej�C�u8��p@P|r�Z����
κ�&�~�.S*!J����
��� �蓅#/s5� �]s�ʉ���	�&�� S���l���
���?����û���b�;	L��'1_Ù#�\8�]l
|YZg�36H�Vs��`_�圕N$r�?e�)>�SU�^��H6�ކ�?c�%t�T@��ʒ���V3�w�x�Ji׍1 ]��f� ��^(�Jv �����*:�uV_�*)J)�D)�1��F�0���
*{Z�>� ��Qb���Q�V�q�ɞ���LP�êYjU�/����GTv��T����A�#9�]�������Dn�����%T][Ӭ~"��Z
m:�,Op ���1g�R��`5N�Ɇx�f��a9�؉�7��ir��<�����f�,%hb�\H��dQa�D��2!����*4�gxx���uC�m�`42^L�\�����_��l%K�� ��r�ծ�����0�I�b��������i������IqOn�h/7�����	L�ר��3�X�wI�Z�W��CS�ߝ����	�
����1͓�*G�:cׁ�3��c�����)�)����� �\�T�<@�"���$���SF ]�bysJǹ!�)���QX����A����bX����rJr�f�BV,>��Ғ�Qq(�Pu�r�t�K�	P�GJ��Gfa�\�6���e��u��5��օ��\?�������ܾ$.v�URbVՠ�V�jzc<��:�� �L4|~8y+���r��ZoF_#&��
�b�����{�#r� �?Z�G�=߳�+Q-�bJ�����n_�qB�3%��,��R:�����O��(�'��D�VLJ�[^��r4H�̓'{(�%�5H�w��Nx�
PM�+��_n�-'�m_��A]1�ޔ�jK�� ���}_>۽�x&f�1��Ę�J3��}�J`��4����o�p��q�~K��Aӹ�X
�. � U�d��($3�{�,V�?W߳�u�$,�6�Q���j�|��5aP��ōV7�sǲr7�ǄGk��=���\x��;B�\ξ]!ħv?jTUcA����]�.�R��?�B�I�U��Sm=�z�I�*�0������Z50��yN,+�̬���z��
��=�|�rf���ƿ��k?�`KN��֩�&c[������}�o97��Vv��ߴd[�Ug?3��ҝ߯1����.{���rT���T,�=��CT�ɺ���>���N�Z����qj#�����pL
@٨�a/�L$�J��Yi&*�$4
d��[ I�c���}8���MJ|�5] J�͠��#"���l�J%�΃u�+���xG0�\��p)Z�z�w�-TP���Rχ�z�b�<�n�ǁQ4k8����M�������.�b8�L�����W�G��~Շ�1��S ��{����A�V�T)c��1U`���X��ơ��#��l�ZF��up���M�|�4�@�:fs.�t:�����}���������8�:�L���g��@$�нk��X���z<�L�vNM��+��0E����:���FfB��ф��e�l#A��7�2�a���p��mR$�ds�z��g@�9^�&����\+=,��{v]EH��anޔj(i�j
;����'�����k(�qy���5�z=:U���-��6Ja� +Ʋ���8(�V��� �V%$x��4d��x����r�7h&%7)�8EŔ�7g�x����:2��I).�T��Q���E�l�BQV�J�M�n�"#�̓�	�e�� ����ܫcШ��Ͻ<`�O҇�,��դ�@�_����מ5�5
�����y*�X�\��B��=��b
W^���B�S=�P ������ͬ��سpp�%��`i�Uп�[��4?BŔ��'�¼.�Ǉ�p���hHl��q��\L��" �`+7O�3_�p1$ W���b�xH`�0�J�t���X�`Ew�Mt���c7��/zM�}���=�̞D�=���>��""�we�kb�{(����d�%�S�%�`K�3���C���X�ug�e�s~=��IĖ��G$�i#�ю!ѕ�"a�Y$�M�S�i~�ұ�xU�-�=�M� K��V���������}�DO�m�����Q4�0Mz5q��u����Am�ݔ��V�R[,��2g�&�J���: ��Rg��o*	ę�>���{MGGG��	r�Q�X>�=|V���E��ضr���"tx�6�s��،���Ab�U��/\ ��9���K��|_��]˜%	�
|?i���Lh���V�_���gs'��3�.ZC��K�ͷ�%\����礣,�QAd��lϨq�xJ���\��{�R�c(Ξ��/�x)�lvV[�t���od�V��lm���G�o�,)�M�XQ��S)�A�/4�w�z���ؑ+*�����H�wu�@��pӀp�4;�:���ƎB.�Q���oӑ�e�=b����:{{o�����D�E��m	�۹��k5&�VΚ���ɍp~���`�3%�J�Lv�9���1�=Vq�J9��M�M�}�I�^�C�}T�D%��
ѓS#�nH�P�|��\��?�b�'2�\��27��H����D��B�g$�Q��(�f�3F���	 �q��AL�\f^���b��\ɍ,,��\+�x2���(z�mܼ�	�xB��	' ������P�(Ԁg0�n'��/V���#�/�
}`�\X�O89�}�L��>{L��:������L��b\��/|�+d~��S��Y�� p�>!���m��I����h�����'=�����e.Ǜ7Ocv6��dc ����͗���ǟ���ַ�3���8<�%+ �x�r�Ţ!K�J�|��ilW��YA���E����Z�P�@���G�v	Fansx|�Ʉ�"�S:�µ����⨘���K�!Ѩ2���5�Νج=�����b��6�~?ݵ`�<�����P���U�2�B���R3b�nM}�զ41G��� �λ�X�~t�Pn���RMηM��Ef�����t:&xDř̨zz�Yh$#;[��.gK�����Ԭu �nW3K���p�s�Q����S*�?��aI'�ĥ��U$��h�&���bB�9Y�築�����6�t#Ruk&�H�:hGd_iV,��Q�^юI�O��	���������v�f����6y ���saymR]*
�hG^�؊�ht8�q\̘N�S�O&v-O��l����`#������V��l"����6��y����
�\� `�=�����
�I{���Btcq�}��嚳Q�9TZ̻\���AlG�=��5������Ɇ���ܛhvDّ�)ɞ ��g<euQY��0vs������'�n�ρ{$�p���{Z�(�#d����-��zHٛ�d����}[u�e/[I���[��\�Y�������b�}��d��s�KԴ\W(9Qrg{N��x2���>�A{��y�Mϯ��C�]K_n�u�*ic�r����?e�5{N��6�/���9�h��'��h+�Kl��|��jS'�Z�:{Z�4�Z������%���
���}�>�
p̤ۉ��	���
���,c��>��g����վ?��8Y��A�i�ڪl�J&�~,=���t����乛�2I�4I�ϕl�Bi���u�"M�4��~��ai�ԎE3��X�P	g��$Yݷ�"�XCU�� �����4X0F��q�ךoKxރV��#��ٗ�������D�ߕ=��>����@��<�n�WK�x/�z�ļ��
zE�k�ǁJ����CQ�2����?�k�J�"��\׮8j����9�&�*I�ǔ�F�$r�㛲b��e�@C*=��x� �lgsΓ����� �N��# �g�k����N�,��5�b��d`o�?�o��\ee]$�VWl���(6!f��S��Is�y�ޡ�����
�BI5��u��Ls{x����"*���$����`�����Ӝ�9���=�c��j1*�C ʃ��{,,���/(��d�w"�G�8B�����1;9�Rx��^@!κ�|sV�S�#�ВD`:_����2^ S��n�JB�>|;1�sJ`�wS��`�?.�û�n7;$�0?�ݷ</���(f ��#dT̡� ����-S��~l���܈�f��I<����_�9�q���8F�Y�U�R��t�i��}�<~�7� ~����$���w�j�0)�e%m���z7~0���� �X�TV�AO�7��w.i$��K��CF3��(�.^���&��g����*����E%)1�U�ggL����e�ª)*���Q��h8��F�>�6# eU�P�m�LTrZ��*���g���@��.YJ��P�c	3�:���_݇* ��DR�"���ܪP���˃�G]�^��r�q3��O�| ���9K�:d�E\�z�N��&��x�jQ������:g5:�|���T��0��a_���7�����P9�cj�
��yt�{%��织861�C+�Ő�CƁkv���n�"�����������.�`���4�LYB�/T�5>	�y>_F�7�z�d������!��3H?��\(�i&%\����cJ���"#��N,�g�a����;�\z���Q��^v�X�����M:�-�xa~�q3�Y�T�d��+�x���r듳X��R�P�魚c���b��x!Ix!f���p�[�����M:΍ Y�L�|O�~ӃAtP�0�V)-Ĵ��(���T^2��������{l_��
�x&�������=왛�R�d9���r|�*>~�N�̺�_�
�z�堋����*���왥<�I�I�eEH�ڽ��Lڞ��[��2;3��ׯA����,鈬����*f �z�ݏ��ro� e2W���OJ<��)Vu	6h*�O[RF�JS���)`�.�M߹�IV��Z5�6��z�}�r�$��dX�f<�!h{InVٜU�Zbij���t��m`�&�&cMt��K��Z�K!}Όr4�B�x����[��Z�"���[���R��@�Y@VI�&Ð�+����oBY�[��� #��{��L�S�*7��3	�6F$�kz�� ��q5��� �|��$~��P.�40��\ ��IBIO.��bݴ�@ȋ�j�w�9�Sא|�A�o2[�$����J����>���-@��V��Q���:�H��Y����B��@9�y��_I�C��~����J�R�:y�t�T�/��>��x��� Iu`�Rm,�)$[{/"�ǞQ�w^�	��m�h�3�#4OVj��!�3�s����$��q�Y����br�*׺�.Z��l�҄�bV��gM�I��(��MC�B�)� n�"J�t,�~ ]�5գ�J���TG���bLr��<6�f�i���ڣK�%*�9�Ĩ������:�P@U���xB`��lcz�$�7O)��u���ӧ�o�2�Y(�);��)��L0�ÜR�g��M٣�"���x���19�e6�b~�����x������ƪ�l��f���OL�ʻ�r�)Xܔ�(�56G���ow1;9�����z������K��O�c�:�i=7�������o,"^��W�o��[b���n�J#ZT��o���E�v1� A_Dg����|�İ2�b����<qc���:��N��crx!�ñ��zg�3�<�HR��9_ F�t0l���z�.��;���k�6��Ŋ��L�s�	�� ��~�6�X�~��h���I����PL��嗪h�pC`b��b�J���6j�� HXDtv��v �%Ú	J����!#%w\��8h��<��QDg��X��ח#.�S܏!��p(�61_ ��"���B����iۣ���� ᗸ~}7�++��''1:<������ch1�~�6V�U���%��2F�z8<<J�&��!m��grx���YǠD$��3ɲ0q��/N��y�M!�H��uH�
2�s��=�-������C ��b�u7N���/D�~����S�]������a�H!��^ぐi�F۬��df@��+/z �؆:�T�k��SීӘ^�N`�Zmb|tD`څ� ��$m�V���?��G���������+d11�k	���Z���~�8�o���n �Y����p�*eh��t��d7��g�9BV�\@�5�5��T1�����C��^��s̸�Sf���Z��I��>�L��d;�G@u߸@XB�F"f�ו���h�7��2!&8�I�����Zg2�16m�ù ���<6'����An��ag[�40�9�*��y>N��r����u�_�[������~^���=6K�3���2�4\*�`Yň�s,��+����Ց��	�]���w��- 6&�U+f�m>�\�$.�;J ���1c9�׽�	ۄ����x�g]�0% �lO�^��M�|�����UC4�ڊ�w�Z�H�C�.���G�H��D�ɑnZBh8�������H�?9������!�-�6�R�����*)�	r�y�?��Z~��t�W�sg�H��O�!��?h�)���d������    IDAT��B�/�vCS�b���Q��Ҝ� ��~X��A�U�F�.��u�#�L#��ub�7f�~�&s����ߧ�g���m��+�%�?3p��}����{m����#o�{�DRC��o�.�_帊�� �ѕri���;Uk��5�n�V��?I/c*� +.��y���06̇�}��]Qlآe��C|�[���c�i0T�`�*}ڟlG�d�r�0�\�z%�D�3�H:|߰�ã�Ӄϒ-;�		,y�Z$��2gl�Lw�¹�E �#<[��V���T����<�9)������h>���b�Ί��A+ڛ:�^�.�9�d��)
-l%L`�A��5�����b��*�NV[k��U:�����K �XÕw��x���)�o|`��� �P1E�������*��� ���P���V9;����͘^�����/��x���ĸ2�|NF)>ؕЉq��t��є���O���^|p��w(X,�b4D _�fv#�ٓ���w�q�m�D�"�;f�	n�4"�������u��o�������*ƓcV���DQ��ll	��W�r���q7�v���g>5n�r����/Hx�
�0  r�
^,��b����M����`��o�!����7�p� L0�	�<V�I�cu	�ٓ�2���9�VRZT,W��` �<._ţ����J�G����O��DHSBf�eo *�m�8����x����ʁG�n�m$�#��f�5��������1��1��{s��Rc5�LbC��� xЏ�h��(��nl����x�� �M�V�X3A`^9����=�xѧg����>�;�P�
��L�#��5�p��K���z�f�T8��HB�+L�f$abu3�g��g?5>���ģ���<����x��W�/��=���C�Ã��t�c�D��j�T�}^�����&���3����Nֹt�'C��L;�q��WW�3����r�����t�W�Ѽ�lr|�+Ǭ�R&��P�ٳ?l�b�L��'/��������4��*���E�	>��4�7O9����b_$�FB�ç���dLկ��9�Zo�~�b;[DLG����'N�,����Tu6km��*�g��A%qj��$�
���pR$���Z1)�R?'�Kٔ�v���AW.�ʬ�������:)�r�i&D�zV�� hVN�L}[���)ql3R��Ź*����`�D&o�ݸ7I��y	R2i���dO�r,�LO���L	^�T�J��JY!4`���/�n5yT�qr��T�a�^x�����WG`?w��4�vy-S���p(\��tM���L"�#���ZD`�?��"B��/��<���k�w�����"X!%ҌE�H�J����T�=S�R��ф�)W��9ŵ���-y.�U1W+"h;�u�}F����(�}/	^��$��=� '3&��ܦT�$'�q��aN����i�
�G�%	;�%�#��;I���z4��/��_�_WY�`�\���/�	���/�T5��|:~8��3tU�ϳ��zf���wl�C�-{���v�kϋ�����Q`e�i���5_@��J$����:#�̵��а����$=�J���:`v��J{���tJ�҂�%Ux!R
9#�:;�� К��3�w(,�\g&r�%?�����g��p8���~9��ָ�K1�ȱ�S����~�$n���t����E,V�/P(c��b 
�8&{�5�*F[
N�$��3 FP��9�ļ\je���̽�Rzƴ4b�[/�P[m�޿��)��@��K� 0�Z�/�#� �����S'�!`z4�j
s��k7��˶B�=�g�8���P�J�Ϭ` &`�׷X���,�(�@)���G S�/����ڇ=��Z~)I ���0��`\L�vs��e��u�1}٫
0����n�� G�h6!P���i,�Ncqz#}�����O�>�8$a��9��I��J�0��t�W�:������~4���{�F|��~:^����r��$%���6�؜=_�y�_�e�W�Id�ր�c�j��v����u�_��`��K1���>����lqLIJI'�4:B0<�q����4��0�图:���'���^�ڮT�I.�L��{����2O�g�5��}s�v��Zڛ�)P
��ӣ���!�U6�!�J&�_����8�YL�x�c.ǧ}����~�S�Q�_R���8r�̦Yn8&���H/7��~�����=�׾1���d�[2a��/6TLs�+;�%��]N�9ϼ'��̧�-��;���@ʞa5�w�T<q0\ �a��w��}ǻ�?~ӻ�o���gq0�x읗�O|t�u�e~��|���/���/P2x�p��~%v�M�.�����~��m�. �*�8ϔD�e���]���ҁx�`I�쩒������Y��wŧ?�)�?>��;�����A�^χN"���_x�ş��?�nt{tGc�[� =ά��(#6%r �H6�3�N#%4850�m9�-t 0?��fH�asN	|�Y�H`�ٱ��������\8"0EŔ3B�r&�$";1��4`�K���|:%	1�p���NLq0 )#D��$� ��U��77Nb G`|.�|�8�(SFutԣ��f��ֽ��7S������g��e�Ԭ���ڛ��]�c)J�(_�� W���T>���@���Ж}ؙ�
�Fa���d)g�ᙓ�F���hyb���t"�ދSVs�j,@M�qO�y~ɹ!��NPs�6`�&90�I���>�"�\MR�8Y���\r�f�?���(kޛ�Z��$��;���~�]7K�[�˧_	�a�M�u��$�6fke�������.Uy�{0�v����I��T���9�q��s��[Q����@U0©B(��5��g�-�I3�[vR����^�M�J	�a��9�ut��і��.+���G
x�I_-)����L�tke�
��譐ץ=\gs��ߴ��<g8{\g�ߎ��to%��G�GM�oA�Ḑ[��D��J�[J���vSL��W��[w\�/��Ym�=wY�zNcM���a��,s�c���]�=��%��p���o�Z�XQV���3�������W��C����	��t5�������*��f� �4�ǚ�O���&J�J;�*m�B��<��Z��K�~>6�_H��Jg+�/j��s*�b�g��9�������5�l�&�`FNx+�;����3`������zy#�1�KG��'��}k<�qw��w�w�z9��@��u�{n����t�g�z�4x�z�����_���x��7��<�7���a�7(��@�'�/n[�aj��)�u��	��<?�,0�c4�8�sAN�c��"��ן�<��4�S;�j��el�s�[�$��NX�B��x�A�zЮ
D�W���"���8��������8=9����A?�1�~W#��ȄkD{r5|�W�Y�`������7�R,O�4���i����dl30ݜ�pq5�v� ~�� �5jP����M0?zU<���d��Yc%"�)wҲ:����$�ӓX�^�'�6����/�O{�c	Lѣ���}}��G?6��θ�	�B����㻾;��̧�w}�7Ƹ�%Ћ�����_��z��c�=�K�pV(�:*{�-�|��7~ݗ�W|�'���$ŷ�-u q�S��e�>g���~������x�����a�n��R ����
V͋e�p�:�g?�	�}�翏G�� �v��(�K��>�g�xs�G�|����������~ ,*����8���Yj�����i��2@���i�;�YV�"�]��Ɠ[����u|�G?>�\�Cv���� [��Y��~����D��P�����+�b�@_��}�j��I#�P �����Q�L�k�����8����D��`Y��A"����7T������_��o�{����;�K��Y������������e�浯�?~���?_�o>;>��>!�������_~]���:V���vG���Q���kc��@�Е,2�;���j)��z=$ޜĝv�_��x�'=).B� 9��]O��7��x�"~�e��W�vx9�4p��L�^s���U�m$:�D��+�au�`� "i~���9[������cN��8�w�g����)����PS KWLӈ��(�> ��~b7�gL� �L7}���4 �N��8� �n����)犁XSK)'XO<�~t/L"$�e�)�g1R
� �Nt���]t��؞-��_g�wܳ�f>��6i���I$wLⳒ@�|�L<˨�ʸ�=�NpLB��Ԓ�ZR��$�ș4�O�ڽL���S�lD��I�.�V�`� �&eU���ϧM8ur�yS&L��N0�,��J�kE��U(pS�q���<�r_B�}�	?+�2��#�t5G�ќ��h��n�~���T-K�/v�M��>�2���H	m��5aS$J>ٛ�d>��(�X���J&�"�r]e�����i�>�<���:��H��J�����K�V
n �7�緪L��!(�wA��#:\���7�o4,rU�I%�����ZJ �H�?Hed���2Ts &��
��)�_3�������@�����hMYQłKѸ����3$w����PA�<�J��6�\kOdz�B�5��h�| �p�/(|�B�e�M���8�x�6!��`��8} ��W�*C�LZ�����U�a�3W��%�U�lP��)����۪����*�$���5�r5�n���6����h�)���]�AV�y�!3��/��<�����kqιd�������͖�ar�V+�%)�&'�?��7�y5@�|_����C��f{�޷ƚ�ފ�SّC)
��0��X���m�1�E\>��=O�+>�>&��G��Gq4	*$AλMЄ�CY!D��l"����C���w�Ge�������{1=�i?��W�:3TW�G�� Q�\�+έ��VsN9Y Ƙn�a%��g
���@���PȘ��tA���(A�#��!ƽ�n����+`�1��L5���*�+�eP3���w0��������717�`�<;#�uŴs0fŔm���I��I3F��b�b���=���1h?,0�+���?���rg���Ӣ���ĒSF����G볓xܕ~����%��}r�R��^��x���J��ø����+���[n�|�K�7_���ş�Y��뿋1;@:�Ap���|k,6��p�"�r>cI��A�C�������z+���Un7M��, ����{���'�M������O����E/U�,��3�c�������o��/��1�1+��Z�!��zZW�P�g�cJ:� ������{K,��8&E} ��������g2Vfm��4t�hk�݃��q^mg�ٜĿ�������A~�� i�\@QU��v%�`9�E�⯽9~�_�%5���	$���&Ӳ�a=��x��n���毉'=f@ ��/�b^P橕���7�������"��{�k�����KG��������/��x�� �T�{�D<|=�5���x�;�_��ύ{�|�6�E����?�s�������Ӂ�w@dn�l0��(������E��ڀ�?0���z�}K/����e<�hM�%I�t��  [)�:���~ �{~�W�O�~_l��b��܋sY�� ��נhτR�t��ZFb+`�+SHj��f��OJA3����?��4?�F^���G���Vf�:9���Ncsz�ٜ*���T6� �H.�gM� �6Iy��� ����R>K�ĺ	Lѹ k����6�ȁ�3�_z���)]yLQA��8IKy,��g'��$��Hа/�Z��܉S]2�ߚwX�s�B��4�I֛�oB�iF�d��ٙղ�X�mu��<��Lq�jn'�%Hڸ�Y������-M��ђ'Kh������ �:�"�J�vR��4U	=���I��4��`O��J`���^G���J?k3VL�̗W���j'�z��G-+�N������+s��m錈š���Ǐ���<�Z3Q~ZxNd�J2��&	/`�Y��Oiأ�T�koH^])X[�V�2�+N��d��ՈdH�9e_$��2�h�S^��P��(��(n��������"V�i�0ڌ� ��V鑠���UN�9�Y�����]9�;o;�[.ĕ[/��]�Ǉqt8��(�{D-����'K`�jU��� �8����V���7�[��R�
7nL���i<���x����>p-V+$�
G��88Ƴ?�#��ĸx�B�����-o{w������G`��)(����y����	�_-׬Ȳ�L1��,�J�jΕ��J�N�zM"R����.@�7��$d���k!ȵ1�2e�J�Nl�X��0�K�3��z����א1�ya̾���Q
AfO�܃ޛ���Q~����6Q���3���d�,"�?�7Jg��Až�y�;~��ql�u:��Mi� �Mb����x��m�QO��}���w1�'0�����R��gH�M�yq�.Q�d����wO�w�����?����Y,��Xla�
�h7ap�]O�&y�������Ï1^n�a������s��J���':1@��r��*��9ʾ�a������L8�c��A�j²ߗ2?:M��=�������v8.�<��dH`���|��&�!��>��:�ks6'�6(�E��#�2������M�L��l�Oc��q���ɷ>0������^��� ̏6p~�����ڢ�TLnbvz󓛱���c.�㛿��_�S�( "#nn��7�-~��~=�{��Y�|F|�G<=^��Wǃ��}��o��x�'?��R�������;c:��} �afi��(�1��w}���g}�G�摊ǰ�DO,��$�`so��j`n(���6�~�m�_^�S�7wt;��t�8<<TŠ�/�9��vC���ɟ�Q����Uq�Gl����Ć2w�#L+37a`���Mď�����~�uq6��Lp�̆��}�Y��;�+i4� ���̐�P�]���)z8���<7���~\:�셎[=+�Vղz����	����V�3����o�����E���Y���E��a�\.x�LF ���G<����o��x������g��	���n�0�����uķ~��į���>�w�|��Ƴ�~E�h�U�1��YgS�"-��1���������?��q�;1��PF��b�?ɥ�|n�a�^'�y����]��Eg��ħ?���������Hy��E_��?B2�QP?��_��E/��x�{nƪwĪ)�z�����Q���b&5��\�n�,���Y1e�)F?]<f���׋�Ť�y�4�C�����5��.��`9��ш�xL��J�qm����8�k~6S���(&�\���X-e�6LV"�,���`:0�˫���'Q���az`��b`��%d{`3�?$�����\��`�'wnٲˢ��:{z�H�2��zP9P�M�a�Z����,8%s��^�*��������$M����'P�{?R�s���}�5!�L;%���8H;z�{Jr�%v��lGc���ؒ�r/Lʽ����z7D>��#?��v���#0��������}���H�ee�ϣ����,�تy�O#��|4��ª\�$2+���bS��{��>�q���2S��&l���S�/(�g>K�6�ַT�����
��YO���L|�$�>� @�稵"�W�dUq爵�ܣ�D+����~�C�	Q���C�wQ=���=ֱ��QQ�^̣s�9z�΢�؈�N��"	ñ|0������ �����A��ʕ���xr<�Iwƅ�^��y��lwl�e_�`�<��_��׿מ��x������7nF�����o����M��x��k2�m�>���_����BiC����?�/^�������u@D�j�Cz1 ���ޅ�Z�f��>*�C���S    IDAT���: ���x����\I�6�&�#C* I���:������O)1��� #@ܿH׳Z�%�`��k͊d���i�����"������Y�R����Ės��UO׽��+�{�*�=`��F1"�#�t��NH������6.dNH�d�o�@���_�ތk ��o�%�7����Ӹ�(��?����g�G=�JAq��� \����[r�Lk)��~��v"N����F�џ�=����*���I�;��9�%�r�^��S%a"�g/"I6C�p��)u��^:�WF�����0�r����^�f�7�BCJTL�)`��y7��>���I*5���ܮ?$`���+���qt'��OF�(4d��Z��cڛ�b=���H�i�=< @�[p���Q#&r�ҐP �x��>�q�����
��������`|��^-G1�B3��^$��3X�!��!xh�U,1�az3�7�<�3��?�c�bȫXw����M|�����7����Q<��;�_}�s�?�Y��.������/��x����Y�sE�V�E n�;gq�9������O}�=tu�»z&B�ވ�'Ә�`�v�¥�|�R\�x!._��HZ�ø~�����W�O��+��ߌ��8n�|���4���+�'�~��^�,n�܏��쏏��ό��u[\�tL���2&�bG��[Y7
^��am"^�S?񳯎�v�ΐ�"=�k�j��}O�D����A����֦K<7�X.f?2�b9(�������P/�ge�m� ���Y}r�D���ϲ��6��������W�^������$F����7�b�H\��l6�~w�E�}�A|��Y���������S F0	 9���Z`[�ǘi��
�;?��������zCtw���O�g���A�U-)�,ǡHO���$��O�����;�b��}G4[�L|?�rf�'�B��r�HcK�����HgW�p�P������9��ؘ$�B�L���W�^U �xh�_����_{c��.D�J.�<�S��i�P%�Ψ�<xdL�D�<0��\:��hL �$0MW;f��c�����k7�����)Ž�����z�u�Ӂ<�f|8؝-bu����{�cr�zL{�X���TD��	L!�tbu�4ↀ)�( �eo��a��0�ގä���I�U���p<L	�|�Ŏ@�&'	.�@A<e���3��^��!qV����<M$Gڰ?-���Z��Lef&����ݛ���
L櫹�F�h��xq�`�V��U�X�!�â���'-Iw=�d�dD�0WQjuHIl�ͪKִ�$#)1�{���4?�3s���D�w&#���U��x^0�`җ���߆!׳���q�b�?�t�˞�Lvy]����I�2���$�Ub�Rm�;V+��x���a&N�o�!1T!u� +X�k��,�
����?ڐ,��+�L0��0%��}�#Ks9^F��d�hL�!�C��<�oH,�8^nzrJ�s�^����ZLc4������u\8���3�\��^��/��9���`�G�a���͘�ÿx�@����/�S�I�j�Z��|�>3ec{�+k�B��MS��+�m�0`Ee�ᇷ�����tL����;�K����r:�xÛ���1�&`������XsuU�MwC7MO��� ""q�8!�р(�511�O�8d0q���A��ST�Zf����z���������~�9ը����y��}ڦ���=�����^{��6�=�GOLa��#8><�rMg*�*B
�14�%J���̊3*�0/J�ӈ'x~�\0�F.6z�+Ӌqb\���<�ޝe��ܾ�B��D��+��gZ�r{ީI��llp���jf��F����6�Z<�	W�	/sp��;��rV�=oA*������,~[H�}h�+�Yl�<W��N���V���3l	��n}�A��>�2�C�}��X$��Zu�,�|A����p�K�aV��I�b���B�w��B�˓�=���xL�-;��������G0Y���a]FT&��s��5��g��`9{�9Z)��.IqΥ��32y�Fb+�ڳg���&�T�Q>��3S���F4Z�v�����+T���&�H�p	J�Ǵ�Fnb
�\ޔ2�S#֙��z����T2џ��8��'J�BW^zz�i�1%P�!�T3?R5&����B>oJyHT�@`���`�ئ|Հi��vXMdj%G����h�	��
�Z���2�>��+��}׽��#��3W~p�:���GQ��Q)��W^����x�����~�_=u_��]�ȑv�"����P-�@m
�h	_��p��˼8t�}�������!_����(���&�E���:�D��gap`6fb���hGX���X��FLM�	ő����rV��!b�8���	�\�B�8�ri�h�X�h�T�����ݍ8�I�O�P(����SOO'��.�ex��P��`0Υl߽�	�N�(�)a� S�r(@pzǎx	�V(0�C;�(����+,U�]E4\C�2����2|��o��Ԙ���	�~ǝسw��QĠB�McX���9hL ���`�D����)�MU���&��E��ҵ��@�x��9��ԧ��pѹg��+��&�
�������~v�;�BEx:$c1tww���s����_��k��萆@�������g���+�����^��
 !�~j�v�O�p�<�\����i�y��0�!|�ޭ����F��V�d�TJ�c�ܛ�ϓ��3�D���3��^ h��QB���4�Ӻ��֗o����n�ۭ��M�oU~+ǣ4���#Ϝ�W��~��G�t�ac���17d���f��3X���W��K5@V�2I��dc>��H���7ނӉ)�ӖbMG�.���7C��t����v�:(s!0-�r�X6�DO�؟�CM�є`�,��ݩE�V$�<�<`��)�/
& &GR�H�������B��8V%{bES�qP��q1a�Ե�[k�f�6dn�r?�,9��#��|�B��G�a�UНR�I5)����N���;��H^�Rys��r���*4w��:7F#�8p��R��XZٶ�J�qC�)���:0d�N*��������5=5�q}��w��I�f��%�~�biN��:�L��(����"�jJ�h��K_=F�wtu�W���"�����{J�f�Cj�VL
0��^_K\<��+(�s��/s�U����|��s˶����=g�+�Y�`�E)l��J`y�j �/f,L���aL����"��a�I	PcC�x�^���s�m�Y��V)�Qe�T�w��:����$�z��`� �.��E�h� �{;�ՙ�f�kˤ��mK��T���0�>�ז4�5c�g�L����f���)��{���� �9fФݮ�`�/}�B�$�%�5�����6P��
02���x�E�*�OL��ɓ:�C�ar�(k�֛<��G�Z`Gc�� ��-��ҝ�H�Sj�'ry=O䞘�������M�=�R�7�[UGX� U�l�}H{]�6��c:�����b5@*�K�X������tȚr'��Ӭ��
���,o?���0�NΖ�y���Jq�a7Kվ����g3	��2�4��m�_�*���ʝ��xԈ{M���n���W��o��熑$�.j9��< ��DA(>�!��i^�j�����|/�\X�x��iᗏ>�{x�Z�����Ɯ�U�E���$n�!'�̃��%�2i���zD����������m�Y�mc*����T���V���1���}OH�����R%�o��M$�%v1`JƔ���o���l��zgp��#/���W���/��*K[$�b��Q5�y_�Gkː��2.��`:'�o|�=8c@[�~K�)�aaL��/=��V�ɸ��:ɉ[2�eI�[(��(oՑDg/[�w��*,[<]]ai>�����>���2��:���<\w�k�x>Y`"�ƾ�Q���q����~��6A�T���H}
�����7��NW�k ����!�a��E������7��G�t.'L�PfϞ��b��������$��8|�"�$�0���%�I�`p�,��:=���j���*�q�-��k�}��q::;;Ŷ���X��v��Q���v��$������_�/d3d�t�:�����j�Rʘ�6ה= Bk�l�h>�S�+�l���D��I�惮�h�3Jk����&�/�����1R��N�����o8zlX��|>'ϠX�������f>a�i�3d�Otc��@;���d^��/�{�EE��ٵ*ڭ2��<��@O����\��k�q�5P�����mx��'�Գ�p��q��O�V�IL��H��w�����՛�``��>��;��c�#���W�����u�ׯ�=��u�˝��ow����wb��nѽ�>ȬP �v������B�M�4ꛢI�c �g�K�,������14�(d%�QE�^A�1��v��O݀���N�h잝�rZ����'�n����b��
"�^�l��fG����Z��d�G��$���eQ�Yٮ�"F&7�)/��{,9���4q�����4J��b?�^������*0�5qԵDV�+$M���t�[L�ʘ&{{�)�).uM�e��0�1�\q��h�Иʣ�zLe��
N
%���-�,T]y�u�A���+�6,��a�yd-������:Aޞ��c�y�j�yy�k�CL<dN��y�j�$�f�ycO4W���.!uL�K�絬8�Ѩ�����v�~��z�y��.�0��s�$�K��:=����#KqWt�/Խ����)0u쇲���LeU��n�)8%y�� �
F�W�:�����;[Eb�f.on�mx1@2��9���;6W?�(,9�{�=���0�Kuu5��3Gr��7n�T��lś��R'�V�~���hcX:��:�%x~������CЄQ�����V�� k��*�B��H��\�OF�0)�ˈ	�n5Q)�E�[)Q�P��fUFM$�m��d08؋%��Ǚ˗b�i0w� f�u���y�J+�%�n��c�SI�:x��4Bޫ���-"���k]����{��6�I}Q;��3h/����������ဘ+$��|4�՛r�k�"��7�Om%���MB�@&����I�?p�������$�G����'����F�o$ӳY�CK&���W������;�z�u��?6�Wz4]\��S����@7�fo���A\��=�?@O�kg�ʂ�'y����e$A���&qϙ?��Z�����
������]`�9��wV��╪�t�Ⱦ���v���"���Sv�����@ټ$��
��*�uN׸7��՘ק;H��|�H3��c���
\�s��|
�`p��?.>�O��2Y �h=~�n�D�A;�E#G�a4C%�՞�	"̹�+�,i4	�d�R��T�U�aK»�T���(N�H�Hzh�5��$W��Dޛd��D������1�w��#�@��4��3���%�jp��"����e����b�^\y�Rpך2_�^(�s#�Q���������IIX2��� �\�xe+�$�Ϳ��ϊ�.`ڐ!,"��<���z?�I���@Z��aJy�*�Q��UnY)�&F��9~$����=X�`s�Q���s�:|�}�2
c��g�9�;�/���Q��3�c#%��B"���D�`1A+���՜FW���}�����:*�@�������Ĭ�>y�$v�އ���HS��+Wa��9l[�6N����~�#C�DrK) YJI�Mtf���������߃F��j��ѱ���A(��tnK/�-�|^dê�
�Pna�����_~���Ҩ���7�����um�=&0��=�����"��FMB�-ý�!�R��(ׯ�d.�	�OK��Ajs�����D>�v��$������\E������s�:�m�C�q2�!���];��c�b�sϚ�C�xB�r�:���3�zGOL�� *U�?�����O�b�dH��j�$y��5�x�ykp�>���N��f�d3��Sؼ}]�<x��8A�_��Օ�uo}>���0e��m�p���X��V��!\r�2|�3�c�0+�v�=���'(�Kxݫ^�?~�kП��C�- ��]�q����C��@(���l��h)��_ho�cu��6�F�c(]��=�fE�<�����-��zh�e���u�K��C�O��G�PHL�v��o���M"�� ˃I�&Q"IH9` �z��}�uRJ�nI��ܵ�N�LL��a�?L�,G��ry�0��
G$	��u!d�Tfv���He�vM��\G�2*�*J-�4�do� SJy2r�=��6k�z4H��hL�К�!ѤS���:R��ĴǴ�k
ӰJy�Hg@��_x�
��c8��[����>��W�Ţْ,j�/UU.'{F��x�BjKd��g����%��ˢ�7M�%	�=����Ɂ?{�u�%~b�a������?:GY?ys�%{�므�%~��볳�F���hL-F	�o�g��s	�~F�N�����z���e2O�of_��,�S5�?�%�.q� �I�����ğ�Kx�0z�4�����J���K��p��Xz��@��H}A6b&3�WL�]bm��C�3��V�q,v��¬�������;lf�$�+�+�Z�U�?���"*�i�Ƒ�x���:�e����s�t�̞݇��[��Q_�$,������p-�~2���,�u��R';��{1C�kx�旿�epK�X�ɳ���pq�Y� �e�|���cx�QAZy�m3K���`��8����a��a��8x�8v�܏#ǆ1�1^,]Q�F����"�4�l�I2L#O"����W���I�ݨ"���?�3��}�b���]����}�-�GX����)E|5("a!�_'�ݬ�9�j��Jm�P���F���������W�a�9�����W�O�We�����3��b�����<�V�����P�%A��S�f���Y�"��u(#ў���Go|�ΏJK�g垓�L�A[װ��ͨ�8�.��o��1ZNB�n��:�XH��_�[��}GF
(4㨇S(�������R#/צ%E)���c�Ėε������$X�U�g����V1ֱ�N�-��F�����9�*0Lt�'��cJ��8��f���TJ��՗��H��_��4?RW^�1u�9+>A�zL�1-���$�1e>AƔ�K1�(��@c��L�baCb��Ld^_C�QD�<�UsS�ӥ�0��o��1|�����E�G�n��GI/�FC�C�*�j҇ѬUP-�f?dSgw���If��U�bɂ�"�Ѫ�P.�FTϾ�vَ^�I@&-�(r��+��r
Lo�.<�4�K�����8�u�m��XE�Z����w�EWW7�`f�I;Q,�06:���1	$]����a3�T*eI���zz�qƙ�E��@Q(�g�l|a#}�Qtvt�o��X0"��Q����H��ͷ����؉jo{��/��cȦ8�Ӏi��G����S���7*��δ� ����L8����	�o[���J��E��72��}mp�,����!�w��r|䆫�1U�*��s$)	�D�w��/�v�ځ�Q̛7�0�?�����S��,`l<�����:J��R�!Ek|^+��ׁ��W`��EH��r�O���6bt�$>���b�ڕ�ܿV�M��m�r_����s��V��=|��� z�;�1�Q&[���_�w<�~������_� .:o��4�������ݎ���c���z�ո���AP�2�|���ǿ��0��٨��{H9/�5���R�d��Ff�7�c��*�Ӝ�L|�y�hT��5�H4&�rA_�̇�d ���60�&���+D��8�L3�Gj��?�/�@+փ:4,d�9�� ,�,3Cm��}���AV��ŖT�Dĝ���1�`*߮�\���t�霮C�e�Le\��rз��?��hݑ��zC�h�V-We_E3g    IDAT������h�S���kyi�L怩�\��@\���;��!e�JS�KƔnx9��`'�)�rm\L�RC�@Ɣ�:8۱a*AT����{V�|J��������m�"�X�#��J�uZ�Ҋ^
�zH�lv3�T�_��5ٯs�S�@�+��|�B�a�N�g3se�C�!)��Ur1IRY������D9��:&��Ӣ�H�X�r�)$��QصKb�-���i*�֫����mA�`������̕e#��p�%L5Y�Ǯ����ʓ2WnIT�U� �+:�ٖ3�Z\r�7I|Oa�<Ϳ1�n�J�1���X��nx8�_ 
x o%)�N��n4�kAq�ŋ ��-��'�X�d�^G�Ƒmem!*ѨШѪѐ��P���L��:�ꬥ8��3q����?�����N
M0�V$���ݭ�n�cq���42�����;E��W����[FIl�Y�bݭ&�b��t�EW݁}FO�X-�0�O��R�F�3J�O�k���Dm������${#�w��T&7�\���\*���p +��`��!'^�8��|2R�-5��cy�����G�y�<�i��Ke�O��ю5�H2�h<Dؓ�0��D<�DL>��~�y��EM�`��k�3Vҫn1TC}0�g�X+縫��>u;Nװ�cꤼ���][L r[fT�����WA��_�>z�n�-�������,�]�����*&���N����U���V�ۧ_�T�#ɉFmkŻ�����o��ӳS�g�]���Z�u�i�<gTl\��ҙ,x���/��bХV[���k��c������x���j���?!��x��K�Q�?q�晝�#ڙU�^2�VX�ϩ���#�8)��Cq*R���eQ�6�c)s�TR�)ӨJ��^23ـig:##c
�S�\2�𼍆��M'U&S6��d�������Q(	�\y#ٔ�IaH=4��z��$6M4j�]�Ȩ�P��H��hy����KgE��R^�Ƿ�⫷�Õ8J��cq��Y�%I�cJ�W*�d	B+R��2:%M��d���V��X��m%m�J �M�V�	c��ږ��=�%3��(�LH�����D���コ
x���#�H���G`�H$��q�4�.X�@\��SB;�'Q-��Ec1�o��({�̡�e�(�J�D���I_�d'���ˇ�O������?���~��SI�
�*��/|��կufX��w^�Z|��>���F'����Ὓ���������� K�.���9ӈ3�Y5&	��Ӗ2��b�l������=p�%Y�2�<���+�w�
Y� �}�X�>�T2�|���_�G}\���b�ra�yң�
����@8�R;y��IokK�r��?�fQ`�¹���63��6v�ދ��GR5��|�=]�^HV),��#�u|����{�r�h��*�tG�$<�t��*>��w��v��h o��7^�׽�B̟�'#T�޴w��cl۲]6�K��MW�]���G"�{����Hf�
��䳐�Ϥޝjt7U	'+�JT����X0uUX�Z�q�ZB�YE�5�����w������Ken��Y���7`;�F=��{��?���&©>�Z6z���*��=�yU>�c��z���#- ���V�{��S]ycٌT�X��O�i��l�(�Ёx��z�(�T�L�1wd���7I).�!zHH#}[Y>��_�h���|> L�L9p���T�Mb�j�i�{����"�L��`�Ub���Yj"&�z��v�l�س��M���6O�*Tŕ7B5�s4�Ky�,&��jm;6e�z�2�;`�x��@ˎ
7 ���Y�����F��dY�k�ȻA�ʢ9P(Ɩ�y{��5%	���~Y3;y��( ^�j��Lyu"�v)��)E5�Af�3	e��H�=б1)�p���EI�7;UN��XӠ�.�W�k��I�Dm��o U��$t&#4ɪw\��%�A�6�Y��b��c)���
,�����<o^R鿪�^.�2(���I�})�c�\�­7�|�?��hK�J��=����3�1��໙���[R̹�5*i�(��*H#Q-!�n�#CW
�g�a��>���b��~�:k���E_ot4gۂ������k'�v[?�٬q����t�����7��� /*��|�̂,{�ʕ
%�&r�&'s8v�$6��{�B�Z��+�Xk��K5���J�Y��d��X�9��S��`�`?�^�+W,G��d�Jđ���|�ӱ�9Y\�����6غ���$�|h�
o����}���V�|Mp���*u�J���<�mߋ}����ѓ��ax,��b�:�q�R�QDI9CR�Q��6�8��������lM]��n�+��nj��O�OT���q��/�8�EG_mq)PL�b�1lԺM������p�,����{j�{5Vظ,W��������~�sƙCi?�[�f�耭*]�N��Uj�~:�?�rv0��z�p��$.\���j�]ޅ��{t�]�3*�3��M.�)���739o����x7D8����Ǟ���l���2ڱ,��-�jd�61�����B��v���^L����l���q���Ơ�cTzL�:�j�� kZ/�P)�dl�54�f!�;+3SY@�v*�:�2��i:%���ITl�$3ږ�{8��)S1@g_���V*�.�PC-_O��2�9� �)�qYX>�1�B<���S�ESF�U`�r^���X:�;���(�n S���q40{GLQi�ې�'�����kR��jh���ё���5�pp� {�j��'�E�X��,�s�j�w�$6�<�[�TW�f2�D��j�v�f}�:����kx�bb�=*&G�}�4Y`��E�;o�\	�2�\����(N�DF��ۇT6+U�������W*�D�80w�4�Kñ���<�����p��q\{͛����O��e��i�ڷ�Ľ?�b�J��*|���3�[�]?ۆ[�z �y����_���1�!jL�<jI+�7�V�������Rj�����R�:����+��^�tT�&~�r�
V �������¦�������G*�Y�J�ZhV:pS�9������B\� �Ӟ�M9 ;:��$谨i�stlw�q'�X�>���]d=.,O���I���G�ك�F�T0`�j|�=oCo��xa����U���܉�7�&�?;ov�����ٽ��#صo��ً��qp=&Rq,X0KO_��������8�#�E�c���^�T��K�fe(���fi�k#�Hj�w4�U�;AXUdu�|_��͸��YZQ�@M)�27RB�'�������O�o��3L5:Ќv���F:6�㟴��p�0gE��֧������Xãn��{Lc�+�����N�l�&P�P��&��h AuCObٴqK��x��E�9�֊
Lk������8�q3YJyɀیU��BLL��h�l��.�=��q1"�$ڂ��b9<�n��F9/�@	X)���/��0�����+-��e�E�#��F�%�Q��,��F�l�M��%�vO�����dI��	�6�W��{�A��t}�.Q�WK����3��SN�����G�$�z�~�4��uH6h[��9��A��7�&ﺄ1� �v���[��l��t�-J�|.[�z�fT�"/�۴����I�]00�\�7�c+)R (Kz`{-5��K�`5����⪎��T3=
����н������JY� ���Op��s�M��3s� �RnM+z�(��"��HGY�F��)���JI�Di�Uљ
c��^,;mV��������j&M�-�N���G��BR	�\����z�%�>���u�E�d�*5 W ��&0t�$N�N!_�b:_B��e�ŲL(�i��Ucm�̵�爎����n+Q�w��G׆1b6H܅�%����#T"I���3ш��!`�sf.�9���LJб7itfS�̤��ۅ�,g�&��݅��N1v�fRl�g�N�g��Gv׭�kg����1�V���Ȉ,eY�(ӯn��!��}�v��-q���5��B�4��b���N�;�d4Z$EH�ԛ�
VI��\{��,���يrE �X&Yu�����ܗ����g�I�U�bA�!mer�U���e�k�׬*8����X����>wu{� ��U 칽o�J0^{�8�Z�2P�������L�!�T2T���e}���ހ��@�#�D�������b����I��{N}=�Z���b����|�����Gp��4�(NN�0��ّB���������S@ϋ�����R��/TXJ+�X�'--�y�H���jy��AƔ^*�0��� TK�N͐�M����R��FM��&Q+V��dO�fi̤��2�}�̷̕7����)s5�\���M�����0͠����b�j#	�	��\h�U+#�(!R����i|�37����i~��u����[�1�+o��bء�eT�4a� �ZBDܮ"kb�~����Rɇ��Q��pzxuf3X��,�w�Jtup�-����������H���Xdť����L?�Q��ƀ�Hf�C���`g��A�`bb{v��Y+��ջ@J�*%�?��ĔP���	����L.�u�v��K���9�� 2�R=�1<�����7��w��կ>~�G1��W���n��v�C��/C�XE1?�?|����G�#޸aL������0&
!�C	��e�@�hq��R��R<|��qKp���r�3
(}
5�������k�����%��oNW�:&���];�W]��[�E
k��f�j�v�F>�ì�9�3o.�t[m�eݐu&3�Ò2����ԳW��j����w�~���\û�z��ͭ�M}r��w�7~�P��Up�u������L�c���B]�5�#�jpCdM�h��$J�<r�r7�e�u����+�\���b�H����f�/�d��C:,�$O�#��S��7��!$;У�/2a��[G�2�k^{!�⣯��jrb(��gcE�,L((?�n��u��ͨ�zJu�Q�-o\��zn.�w�ɜ15:�(}�cJ^���R^2�!�PSFL�qfo�������iu:'��ɧ�&qd��ͦЈ�HwH�{|��n�Z�b�\uZ�3�S��w!��S�"�L:���X܆�.sI*	���T�F1�-����7�cG��i�����L,"c!sK�V��P�)�V%1w���Ȉ���@�0��cpS�-���Ur;�Q����Ez(�����S��}��'3 ����Y�04��m�T��&��./��05�$/�w�X\�[���͊�M8��Z�/d��r_����	������_rO�� �k׼�:/��f^�����p#�P�fZ�?��̹в�`�^ e��PV��m���1Lr����{�W^L��p�LV���X�"*�tEL*Z4)��^d-���3|���#鑤�r�z�uT��� �,��ј��[�V����Z�Fyj�
ϩ���8}��1g��k�Z�E���q��z�i��-0{{�T��d�n-gbu\�c<�j�Ɖ�<�'�Qȗ0=]@�TA�XG��N���(��t�Ų����O�!!K�2�ˤ(�"��qo��
��38����I-�����������W�-Vt�Ձ��ǯϷ)�wFS�����u��@<�5R�6���tvf��׃�L�]Y�vu`�yX�tN_<��'y��73�*y.�'���̣�͸ރT��B� �
��)`����y�[������T	�p�x�T'b�.D�D�I��)Df-��-|�X,�SZ�N�	[.�E�e��E��D����s[��On+'�����͎�)y���hy'����p'�TX��%&���b��ea��!�2�k�?�($y��@��3�p�:4����
�v��^���͊�vx�U��� �l�?���kE�q7�'���@�+����R?��oݏ�#9����8ۈ�h6���u!��3��0$�ʸψ#����25z�H��I Z���sʘ�,b�T��d�;g0��!iy�v븘v��eX�)�-��cd�qtq���2gj�Y̦�XX���!�q��2_�e>��E���]���+�Z�:�ś� �p:�P����O浨���TiX��R^imb�B`ڬ ^��Ysi~�,��G�V��E���m*�=YI�܌�AsQ4h���I�PK�k��+=��������;sn�靘�CR�I;�\����<��P!���D`��D���a���j�dtn�8]F����?�r3^�j�0�Mj���ay���~y�j�"�����.8]�ič�i�\��ѣ���2C�� b4>ⵑIRj���"ʵ�v�����]=��z��w��6m��^{>���a��h8����m'����Ǉp�����7]��be($�u��p��~�r����%�=Ⱥ�}oK�M�v�R��s���,g����)אU�
𞷿o}��HQS!�an���5c��K����۰w�n���W✵+�U�UI+��81���7J���ۇY�x6��������PdB:g�<t���R��������7��U�V�O>�,\�@�[�O��XK��/yVzLc�2����߂ެf�&���3_�!��p@^;��3�L
�$C���p��BMP]��(��g���U��Lg0<U��߆�'�ҧ�
��s`xL��r��$&�����!��|��c�Y���*�Vu�F��۸��oĹg�(8e�.j�����1��G��~��|�_~��j�vZ�P,!�+̝s��GwЈSm�f�dC3?��sK�0D��^��)��iJ�RK��^dL��{�p��2��Ŕh*!sLci�YW�R�C+��"I��5Dv_�q܃L�����T�i��Uy�X��ڗ�O���4?j��(�7q�)(�tf`J%DʫA<$�<�R���̐A�@`�`�^�9D�JV[\-}`*�G�nX�^M<<ӱ���J�Ȍ�����Ele]]2�ƻ���@=(�I���TΥ늯�����������7�K+��%H��L2���êy�z��8Y�b�f����s�]w�xA�U�dO*�A�]t����L���:v�}>gH"�ԍ��9��VtH���(�̥�hǤ��49@ȿ�M�T��qM�2��ΙyR���tN�ܯ�T�]���wVt�U>��Ip��3#���1��*�5(+ZiNO}~��r3<ƣq�9�)�'}D�\�\�JS�h��m�1�;) ��sV�����ӗ
����W���-��I�V�ZԠC;�����Z�N������p��q��M`*WD�R���4�&�����g)�E�WoE �$�~'R��R�*U6
��$,q�D1�U�'�6Y�<K�&\����s��c�w��b���m�>ng�Z��$�	���j�^�v�皌yh��u��Z;�����~�;�F:�@&�܁^,�ۏ3�/��K���әBWVG�˶+Ȫ1�5X.P{D�������%`l�����x����3�q�d�J�p�T7B�,b��TqƂ3۵�H;MP%�����y�ѵ�6������"���͐MLa<���6~�w���
H�}�RSm���{�o�����@�)tXҮ�}���u�͟�n�]�+Bz��`���z֪�9�7�n2�,"����5�������ėuj1XH��S��7���������Ňz8xlO��w��cS.�\����߄!�XF(�~*�d�c`:�t_���jҲDܠc픜�\�X&i!�5T���ˣV*j~ߊH�S�3%�L�Tr�6ZCY`�9�%0��zS#�L��Y0��E|e=�o�1���	���e�!�*1�3�S�gɘ�<W~N9�m�R�Ap.#j�x�z�F��V�1���?0}t��b=��v\̏L�$�"7g�$Z�r(�mTA��Fag/���?y�Đ6`\��u��V�4孇�84	|������Pi�_@�躇FA��l��ŏ�ܕ��arc�r16�H    IDAT>!fG]�=�'�O`t�$&�Gq٥���Sf�1�o�8~� JS9�c1��"�e*� /@п�����
��R�#W(0Mg�
@"2M<����ޅM7��W���ǂ�s�Q��ގ��h�ނ��w����x��k���(s3����܃���(Tu�/��8$%�Rŷ>�{Y�~;�`-#bY�)����@ X�X�Ai�px�p��+�$0m+��\)׌]���a�ٵW��W]�
�^��ŀ�&�#G�`�Ï�)Co_�I�T׮�V�J�C&��v�ڳ+3��~������������~�#�W\�fR�����߽��ۀ2�Be��G�ō�F�|�blt��R���HEn�/�+_y�^u���f�<��x"���qU|߮�Ntv�g8|���p�#P��lZ{��mr��2�. �@i�&i!LǔHq�F�ש���5mWs�#���^�w��*�Y�#k�1��0�B*X4j�[�M���N�=ZB43�f���Ye$��`�$�׿�,���D-Mu�UeXlQ`ʠ+��Nm4�����R�FG칠4/G�̊ܛdV{D�1U`��Y��z>7�_�+u��w�>�J-�.]}guI�=�U�R�m��K�L�\�S94ǧ�&Bi-p A
��~�`��Q2!���\�k3Z���q�6kS�� S�K�����.��ڹ!�I��y#2�u�4;�i֏S�00�{�$\�g7�-XĐ�ߊ�iI��V�=��թǺ�uv��bA@��I_SfKج?�3�-�1�͙Ը��Cr
���y_�Ёo�>�z���v#�!����<w?��ս�/�u��K�s�zt�eN�W�eV=V�����3�"�L�I����R���fk���������%��	�ʗ��̱{��|mq*8�EH%���㨚�����H{-	��d���;�l�1x�+��h�j�W*��F��d��x����d~�_�kV.���Aow��*&m��؏��E#rme�i�Ǹ�FJC���/��J8z|��a�}ضc��?gF *���<�Ɏ��w4�pʿ�0��0����Fj(�K���"GYh�GY�L�]��ā3L�|ɷ>��������F����F�{�>y#��LEi���\r2��4�Uɳ�iU�זx�aE��j9�0�h����La��~��z�Y}&��O�+���$Rq�k�^��J`������g���Af{xش}�?�	�v�ɉ2rU�� �Dv��I1N"���9ɞ�*����`QI{����*��t
�ϿF�Z�
��t-�f�bs�3˳��
	��f���G]Ae��F`��>z�LW?����x*��Z�&�V8s9�̚��φ⒬��G�!��5W�W_�n>1�K�t>�{�3���i`�8���6�M;�M��i�<Q�d�`��,�2BF@�$W��F�aT���Qdg�K�P�r^�<Tݣ���$��&���0�y(cq@WF�SǨ��Zy10�	LY��L"L���q5�c��i��4"��]��<��)U 1��!�JƔ��&0x��H+����[�d�Ԩ#�(	0]� #�t�,��u��/�%0��m�����&c�R���b�B~�&�#�m���5DPG�����>v�5��%���唥\\�'�uh���~�{� *Mv߫��i��)� ӿ�^�r�wH� ��ΡP(
(�r��!��Q3�^r!���t�ap�����獤�G��<�Vkr�ku��p)T����L6+#R(�-U�x�Gq�=?���pՕ���̛?[E�YuDq�DO�߉m;�aߞ�좕��7J���w!cz��v�ֻB��D+�F3�F"��`���LI�S�H`��;?e�E�:wJn�	:M�e���HG�Ȅ���o��.[���^5�`Y�Pƣ���g�o�~�غ���R�Y�B@�j���?y�({�!�����F��I�����j�T�"e!� ��3���ŋ��K�Ϭ��~>��[�9��o�u�x;�W��8�4���)Y��B�P7������ף�S�>A���u|�o�į��! �3����G8oM�HIXu���C��b���e�2�LՀ�ܽ?��ch�٫Iy5*������:��#W��o'��V��$�t��B`?G�k(N#Ҝ�9+�u�|	��d5z;�ʳ�;�B ���-���;�'�hv�ΉT��W��+��}�2��Cr����}�ne��c�����	LY���t%cR^��&X(�3����R�Ϟ`�b)��1�k`�dBk����Z�J�����@�8�����T�z+n��2��]=�'��5�k�כs'� q�k��h��#I�
��H�)y�TY���͐��������ȍԴK��T�4(: ��!̚Ht]����'� �RYo�U���\����:����B�`ȀG0��]فK�g0��(��un�/-z�Q��Y��qX����1�� �̐�:ׇg�O9�� 0��\`����)�~#yO+θkU�֗JJ�&�Y{;���9�^��\_������ͳ����K����wL�"n0	����12���f.qС3=��/��,:���5�4�8:'S�T*�C�9��N`+ͮ�c�M�_���bA���RRDOg�W.��.��3`͙�1o0&=�n�hP�d�Ui`�\=R%V�ʘX���Gq��	;��\	Ӆ2��&%ia�Y�?*������,RJ�N-���r�YX���JuR9A��4R��o0sl�g<��]���خ��R�U�zؙޫ�'[wT��f�,n8 �kOG�����y�?P;#!)2��U�[u� ����(�L�f���e��M̟ݏEs�q����?؃�g.Ƃ9����Aa�<g'�u�4�����q{Ų9,<�?\�֝Cظ��}a��Qi%��"��UCj���޶P:l���2�Q�lf�ϩ�T�i�H�;{\qS}��Yj���'ٳ��~�u]q�SK`����m�Y�NН_���s/�ؙo����p���	�"�b�=-��3Y;2"Fe�1Ω�N�'��9�p�5W�5s��$ )n��_�/8�]g���x�7n�H�i8:��s���ɍ��}��s-�*\�)�B,P�i����mL�Tv��z4����2�zȖFDڜ�,�%��2~&ޙA�-F�!c*#c� �R�N�Z��q�Je����ʢLGJ��40b-MFՉ�Xs�t2�$��MM����l���cf�q�9����l��G�Kq�2`Je���&͏Ʊր���0e2GP�Ȗa|���<`�sv�U��_Q��\�MӔ?ivjU�������_�?���M����^��Q,���$qd�)dR�;�$~��&n��xf�Ԛ�`�Oj�Q#cZD�6)Z���8�,���p�I.�G���P����*�.z����dTJ��R���rP2�f:;E����ė�G��J+�J+G�����WX5>��|	?��L�9�k��&|�7a`�W/�����e<��f�=p۶l�k�|	>x�5H��6 D����N|�?D�G��4�[t�ƈ�{Et�̖l9v�FHX�\�U��a�$�?�C�Y��F�i�1������+<���j>��r��=v���`󦍸�q�ڕ:����v�#x��OȢL%�L�����c86��b�30g�|I����� �O>z�8�^|�E�Ї>��Y}R2'cJ��[��3<���(�i��߀�{�:��� v��&>��;��3�%X�]� _������(�&�y��';3�J��& �c���w�{w=�f��h�]bp#2h�����5
� �O��6�Zz�i�ED���K(��k5��L�����l-�Y�=]d��Uك3U {j3���c�yh�� "�Di�"�by�����N���u�"�Qc3��㪚LE��{ܖ�ZqZ�ǩ��f|��. �K�7d�i}:/��\���R�]h��ԕ�}O�w!�����j��N�Qc�<E���)��0%8v�T�	Jv[-de��4Z�ӈ7Zb�$�Zi	�ār/2��xT̏$c�, Le���t��!�n�v�1�RVFÁ���f~dr<I�0�< ���9�:7]�h-)01�`1TVc���=2I�Z> u�)��kFB�^���>x�ϐ��"!���<�3���Vs�8bF[NF��{~z�t&w=��]W?�/Y��2Y>�����7~�K�| !�k�Dje��F"H��3rҊ��k�]Oe`����)x��!����`�����������Ki�D�>Uӭ`V�'T��c*�S)��-�^�gvfY�(���p�d�& l���c��2�Ţ��Fi��*��g�v�b��⳱v�",Yԅ��4e��u��0�^u i�o=k�B�#�804�[���M;q��(&�K���$���=O6@�b�UP*��̙U�'k��&
P��_�GS�� _Lw�\��Xr83(���o݉d�׌(e9z�u�j�#�Gi:�&�V{�N:���5n;)�����,���QZ{]JM9]A���^a~!��:���O^-�Q+�zIr8ԋ������]�W\z!֬:��@)�彔�Ǭ���Z�rc̜3���Ҵ��O���a��!�߲{�F1Y��I�<�M&��	��0�g#}3x��[�p �g���W�S��3SML` >ԑ2ު�wл���]�]�P���XT!/q��y�%c崭�}eE)�~�5�ﳟ�x�?�▎��%ĺs��9q�.,Rp�7��8m0�+/\�����8}^�G��L����J_�z���~�_�s3
$&�*ֱu��ܸ�l>���JUf�)4�1�&"�v+T��0�"a(�]�e6z�T�U�mEԨM�I#���Bu!�7�q1����F;2ʈ=��j#K�d�Z�05�5��;�G5�Q��7��&x��
JS�L���]2����<u3��[�B���9�#Q�H.H�H?�
��1�]�����z,�Z�w0�A`��[��*�8L����Fz���M! �q1j��9�4+�ȏ�'µo�
]p�z�Q,��k�lݲ��O`ttTP�������êUg!���Z�|b7~���>���^I��t �h@7�0���7��I�s���rIc4����$f�V�cx�$J��$��]�T2!��MѮ���C�\D2�772&\Tαp���!3>9�r��y����[�2Y3V]�������ch�>�����w^����9��Bx��������ƻ�}>��w�����v�6��=��b�HJ"3�0e��:�����^���o�� �W�%pr!�*Rь��pu�7��oz)2� ���������'�u�f�{�Z�w�Z�I�38�)�GG�y���?����V17Q�%�uD�N�@8c�r�1�fjEzϮ=��_������W_�n��f�F���C'[��m��Ba�H7�����
Lyo`�����zn'�*�X:����M8m?���7F�q��
��Dk� �k��d�|��q�Ϟ�hG�_�� �^`�e/p�4|.��R� .I��q���0``��6�(�(�P-L�^�B2�D_W
�z�0��+W91���x�Se���F<ۇtGɤ8��~�>EM�hr�{�;��ALp`� �Hy9�4�d�Jyy��׻`LY�`��rD]�&i7��kq��ǔUE��RI刲�t��u3���P�.�b�+�� {L��]y��i:�<'����<�?ulB���Sg����>Y^S����@Ǚ��v����E���)��H�S��3ő���= �
�KS���KAg\I���r@�E�^��}p'��hߓ��[�j9�2��}���&�&C<���n�DJ�ʪ�ueH��͵3�%_��n,��pj߫"@2�Z�VfG�SQ�8p��'Y��/c	%��DO�������2�k���6pݴ�P֘K�g�1فf��.!R �̫�z�/'���4)1�Ԙ:�yqĒ���<P��㞛��[rl�95F��/"K��Z�G��Mnl�i�c�*��Z�J	ਗbAf��tD�dA?�;g.�hV�X��~�Q����LwwK֮�9z�2ӷ%m�(WFjظ� z���/cFJ��K M��=��$�X"!���|�י�{A=�s:O�Q��Y�l6�Ie�)]�?��{� �J/������F�^�H)t���7|`�z�`J@�It�A�}�x�۞�}��-���YWƔ��n���"d˅S�Ȳ���
Զ>U�γ�c�Rh���(�'P΍�Z��d]��.���]p.����t!z��`=��N����[�b #cutip���T2�u W��W�ĳ[�����u`�S)��6�EF�2n&�Y����Ԋ͖�;Way�K:Ձ+�(}��5k�sg��/pX�r&cƞ�Rt���|9���1���xm�*��clG�5hq'�s����+���8��
T*g�K]0e��h�<o��\\~�J�g"2�A�wr��s�
k�_��SO������]$oC'��Ćx~�!���t1�b��Gl�b���Q�E�7��5���i:!��j�P�Z� �
INBW��b��
���0�"��(��A#�SdLI�58j�^<!te��`�R�!76�J�$mG4Cƴ3%R^Np�G�Rd��7C��+2��S2;^}���k��W�	��w�TF�y�,4�2&��xJ�Ѫ V�ً����͘�R��R޿��{1RM0%��M�E#t���	L#�a�`�$��Nc�Q��N�'�isz�l�q­7Bؼ� �mݍR>�F��p,�9sga���8��%�D�(V�xn��8�L�K�X��v!�
�5J�'1���W�kϜ����3���	���I����	�����w��5H����\�QE~r���|��[�������l@��~ ��R
o��p�o،/~�oq��a|��?�7����P]>8�X9���'q�=����#h7���{ހ���Z��ɘ���-��?��ru�e�Ȭ+KHU�aFTL�E�`R��¥�q=�-!4ki�lFn��(>�޷�}�^�sg��|�G�V�� �?�|!��7�g�ܳ�h�\��(yi���a疭�����,��r�.\�\����2Q�!�iK#�Lz�
�\�ֿ�O�/������,�4&�cr-�?Z�?�� |����$�c*�Gc�����N<��vT�EtvFq��^��_�+N���ބ(O�G�prt�RE��s1���D�5`�"������mGKv!a]+�vӕ��*�S����]0��G��Q�cܩ��e*+�"��^A�8�� Ԃ$|<���5�h,�h2�T��L�:�U�E�(	KW�2p�ʻ�fr	�?gտjw�2�-J��ǔ��
L���|��I`����Q%�[W'>Jy�n��OƔI�T��e��C�3ΰ�:_D�ξ2�$:���:�U������S���h�O ^o�!@s$I�����0��$��c�ʍ��Y�*�ZLkb�$��1��v,'�d�:*�zM�P�X�`֯�y�rB�0u&)^_�{D^��?32nެ�@O�K�iΦ HS�NM����I���%A.y�v�&Sz���D鏜0��k�W�3$��m
d�3�L�v�
^��7j�SI�\��zt�s9P��Z�7��X�g9`jW4�r��%ƺ�u �w��'�y����3�=�v���k�L�YK1Z��S5񟗻{A�E�����^�7{�O�q*Z�(O[9����fa���78+����,V��/����z)�Ή�#�ȐIف=�T+X�,���n�I&��gD����0t|DƉ��C'���qqQ�7	c��;���R��~P�P2��>�*�'�,�J��
<�if�M�iʈ(3�QZ��DΦt��Ӯ��
�����˃u�o������g��^u2k={��}�;t?�x���=��v|y�٭en��9�9-@��V�pJL��v���&�"H��Ⱥ]��x��@)?�J1�J)�F9/�+�Dg�~V,_�eKb��YXr�<�u��3&n����AFU;]���J2Y|����I<��fl�v����Ԉ"�@+��bT��rs8RN�j�V�3����%�    IDAT6�n���ɨ����J&��c*U��b�k!��P���/��؋�>c����������a?cq߭[^������]�3U3@��YZ�]��hU�Гn�5���7������Z	�]Yu�����o`�Óe��� ^�y[�ǉ�2��*�j0�1*�dD��F$$=����G�L	Z����ʴvqǘ����VK%eL�Ʉvw �MK�*[����=�(����8�5�R�+LP,:�\��h�3���cQQ�'��d������t��QH�5�[��71kk����%���\/K�i�:�5����h�)m]]�
��P�M�`J)�n��Iy)���Q���bT�C�Q+��I�Q�����I��ꗿ�_r��;q��~���X�a�&&���t�\��+��y"Ó�wb��	�ZI����^zK�E�Ƀn�����Ҏ|����H;�:E6<6>�R��eg����K�(�azl��	1���헛/Zlk��CW+�5� ���d��Y�P/lَ[��ULMN�_�,.��B]�Lfi��n����Gatth���^����R�R������yX\y���$�a:���_z}-�bW��"=�Zю��c����&��f��v��*L?t����^.�T$�U[�9w�\a�(�}�駱p�<�]��X����R�у�pt�X�/[vb��#a���jLf"Qa�;{zՒ�f���'�|
��O�<��}�X�z�������<�~
����&�����w��i�ܔt�8X����X��V�|��������Ua���x?��ظi���9s񊗿�]���l=��Olů�؍�<�<{Kً̽��#�>5�ṙnRw��1 ~��C�fU6�֭aޕ}ŭ�^W��	P˨��r�;�(�-;Dbd R����y�f��y,���*��.�Փ��d� ��TdL4&˦D�KW^q���(K�49��Dq�[0���*� ��)�r��hS�Uʫ�uQ��պөi�UC(*��1�O,�˭:*dMMn&�H饍 �d�i�cL�������$(��@�#�BhP2���͵��Lš[L�(�5`�3�̏|`J)�������Zߩ&P��X\2��i�Q�b�<�@D�V���p_;ilP,�#OX���.!q��:>���H^〞eAS� �l��7�[�P������rɳ�� K�3;�<��H���(2Xkt��;�[$�^+���},�T���1�%q������1N*�:e�b*��؟�F��O�Y�x�/П��2��h"���UA��p�����i6�d�,�˺�U���h1��x��+"�mT�����(O#�,!�b�`.�`%V-[��K�kk__��& ��o�vyl�3�F��k�
�-�89��;�a����8��d�j��&�p"#3y�	H��w���]U���S��LBB
������z	A���X Q��j@_Q1����	i/E �B�33i3�̙9�=���Z{����$����7\�LΜ�<�s߿�����k��	��Z!˾6�E��� ����f�\�\�B<K~�Zg�G9z~}�c�ƶ�c/�3��_���\2�zs���qW�Ԡ�=1��43[7z�6 ]/Fȵ_�cR�L 0-���h����8� �w2cW�g���b�~k�6�m��p����%�m��� ;�Ų�MmԊ8���x��8��c��3N�)'�[����o_D|OkI	xn�F�g/j0t�>��e|�{p��w������I�*�Z*�k(V�� \b!�9��)����-]a(��/��y�(J��=����L�z8&�bw|
?���A$D���	���ܔ��ǽ�A3������b� ��'i�f��k<�0� �e��R�+^x).{�Y�*��u�}�f�9*ɟ���}��ݠ���5`�9����v=�o �=���v�ۗ(��o*3,��@AF�$Q1��V�쫡_4O���-Ĝk9�n�ƒ��l]⸖��c�ƪ�������K�N�p��SbL+�w{X�[и���*n�Ԥ��R�zL�y}80�q�^F�\0]_\0�I,���	��\w)�U���I1@��9��q-�P�[0=���x�o���t��dS3?2�T��do|S����Zxp	�v��Σ�_Ey?���3��7��Y�_>�����|̠Q/�g��\�?G�@��*�/݀O|�:,�Q�3T�́���Ř�8bj����o��S�r��67GI�P���-\��={TI<��cR%%�fg�kV����Q���2�M�C)aZ5ʡ�(h$�;��&�������+'�w^�{���)����ˡ5 �����s_�:�!�U��g/��^�<�m�
�1�����`�M)uUɲ�Ÿa��L/�Imh b���~-�SA@�<�u1겂�D���_����|��z���CI�P�V�
<�V���o߆#vl�5�ßb�FX]Z�=�w�^�ᤓO��1��i���h�Y��
My�<n	U0м���������x9�x�Ė*��>��Z�Ǐ~��ҷ����Fm�׿�x�˟+9��,�]p�{>��_w���x�¶U\�����?	'�t"��w���p�-wx�}��x鋟��O?�J��=�k�z~p�ƹI������\+.�J��,!������v4�{�$��%ِ��E�!�Q/� d*xp����0����ڍʾ%����_��W_:�n�H�!\zk�A�ޤ��=�Fߥ��;�]������f��y�m��+o�������2��Pn0%c�9�T1�P����e&���F;uVLY�̣:5��#6�2��>zyڳ�5�,��~@��0�/��)ͯ�	0U�q1y	P�%$�jU�n>�x�i�]��s�D��^3W�8�N�m��S���n�s�qCv0�y�,$�Iߥ�b��ʊ������Tv�&g|���Wg�<�L]#�8������a`�^����O�
�K0�a?�ɐv������fO��M
\g$�J�#�	F2c��{��_���8X}䁖�<�I*� 6I��Mp��k���91j!�ir�D�^�|q���D'�+^�%�Ζ&�'�d��2�a��{�QM�`�2=��>���rh�-��2��R_������3�r!�:u;��6k�`�C^*OxcB�w}4%�4/���������܉��`a�)��B��+'Q�L _�moC�9���EP�w�9�T�|���~�'p��j&>�Vm3����P�x��ٳ�l�y�fz���K�c��� ���P$ڀ��̈́���:��vU��h��V�U��y���:�Lm��y~E�	6� ��vgix�0�6���I���uřp��Uf]n�3b_�96s��~�u	�� �6O`�t'w.��p��g�c�h�m����evUvy�����*^�uuf�����/_�[�؋f��r}�̒4��P�U(�U����q�N�Sd�\N�v���rS�eYj�{��T�2�5�;�~��P�ߚ�Vh��� ��p*tp@�r��40�o\A �O=�����QX� 7�"?j�0X��;'�_��y,*cKL�j(�o�}?�<�1�C�Z�1xhw�7ݱ����r�+tLi�Ȅ��)/5�@�Fr�oۊ|��a��6(��j_�:L���U�c���8&�-�V���q���K`�>SJyL:0%㺺@�<���j)0e�ҸLM���[��*��J�5���()��uK���
��H/�*�����l��m��6��6��E�s���c���vF��k=t��Y���Œ�^k���Q��q���o��gp��D�r�.��/|�|�C����<&�%�쥗��/~"v�<��|��}	�����`˅���i��4��e9����&�>��Dʫ�@I�Dlk�=th7�t��QG#��u�&��e�����9��5��4A��dL&m���޶eʋ�ّ��{����'q�9gᕯx���y�;��������/���+x�/_��͋�S'�b�~�f|�_���^MR^R��3�z�ǔ��r�88�
�x_ڜc�	V/���.jX�[��2����k�l*�K��
���L�+ǽl�4i}kTEfqgh�ڲZ�m�v+lx��읤d`jj
e�$�8�d�z#\}��8�?����ŲY:�#��$��>�����|��f0=��k�2��g`�͡�c�k�o{����߻S#	�l.�~�E����أ&�}�}����'�v˭(�Fx񋟍_y��q�֢6����k���n؋��&�1�t"S-���p�L괞p���L��[�Mb.�Q5p�>ː{E]��^��(l�P4���7r���H����4�v�=z)yX��7Tr�=��bn �6�9\�"�D��nu]��G��%�?S�3�2>�ѭ�`���1]��iIy''0q�U���1�$=�z4���b����:���p���r9g���_�ĭRưZ�+o��1f*����s0�a�4)�f<{�p�`ʸGj�
Z���o�G�o��\��=��`�#�,`�2g=�?����}=��nw)o8�f��GdF7�����YE=5���e~�ϳ�1I�u� ���?#�05y�F���Z���$�CI�<�� L����Ͳ��ّ�?�O���MF�X�&~ ����5�9Ń��ɧ_~p�)��ƎT�a�+1�I�ap�A�۝O����L�L�5Dl4�)��cLS�NK���kKh�.�Z���u<�'�yϸ�?�x�n��ޣ�3�KU�d�)���ŝ!���{x�9ܽ�~|��7��7ފ6eG9�)(�R�@�1�rm#�|	���qabH0J ��2��K�i���]�wP=�Jڽ�>�y.oHLcb�IЖHX��Q[<Sc?a/r,h'�6�:�TRl�m2	e�#��a f����k���3�j^Ψ��� 3>ȁ��,IN?����g��/�&\�R��Ԕ��;��iIz�sɒ��+��lײ�4���|���G��+f�5��o�FJLO���'��K�t>�>�$�t���<	�2�?cn���B�.�J����fx�1��W�Ƿ���g[8���z��q����k�^�rE�A�LXha�A����32S���_���d��2�E�l\�ƶ��:3�xm��ʖ������HX�ZJ�/��3	뻁���Z�zqc/�
�5%0-�0Qj��7��o|N�9��ft��_����\���~7\�Wp���s�A�;����.Z=Սȓ�R�A#�5)��Gm�IyY�f�C@���2�5&���&�6��=�f�Lk�m��w�#t$�5CFF��zU�G�NW=�d]%���.E�4L����S.��D��F�$u�~���Ӣ��'9�������E��>Ţ�����حk���Ұ�Jo	�?�?{����m�D��RޡKy�����f%�=�)͏T����dA�FjNe>C���2Vf���Û�9x���-.���;�_ſ|�Z|�?��6�qO}�yx��ᜓ�a��F����;���~��쓬X�ƛ����m�Y��My���o�9Y`J7�f���
43�����v������p�M����!v�1������ip�殻wa���h�z:<)/.��@R��%L68ꨣ�e˴)Ӑ��0{� ܷ/~����^�ʰ�߂�(��#�џ�-��3_����doy����S��}�F��ǿ�f�&�#.��r+7�f�����J805G� -���������8{v�D-���y���O?E�\� J\�Xmᓾ-�e}���sϽ	Sc�V�A��t{�Ӝ=4/�+1x���9�8�;H�=��cp��'azzRn�d}��q�]w��>�	<�؝��?��C��1�ul�����������y�*��e��/����(�صw��]E`zƣ..8���Oނ�)k3Pf��/݊�]�!ܷ{r�>���y��_���
����m+x߇����V�/ptG�� zG��X�1+�z���2O �Hz�7P�D��/����,�l�L�V"�ԉ��]����uC�jJ���wN���$)PՋ� �ǴǙ��j��
z<��o��z�G�T�׸������q�2�U�LX�c��0�˱C�� TiP� i���)m�kN40�c�������K��+B`��t��������ס�X�xČ��\yK`CSN)1�a�!��J���]�92����#��W�j������D/�0���¶3u����xOSf\W�u��I�2��#-RJ`JL�Ǟ���w|Ⱥ�`�u8��^/��I���9�{-a�Ҵe2�4.�3��o�S�5{6	����LO� ��M4�&�N`'ʚ�
�۽P� :�1�*]6�F6���P_�5�DZ&�c��+��%���&}��}<�9�?�lÌ'kȤ��L���J.8��������$����.8�\t�cp�1@�G��=C�'���o��ڝ`���{��9�[�?��ܱ��[�`�G�XE�fE�-WQ�6�X�$�̌lTK:o����N�r��m�P�f��uЍ7�T�y�@���PBH� �L�]�sJ$��X.[G�
vJ��YS̇�i�zj�w`�n1&qy3g4������
$�gm@'VrF%�d^��u�,Y�����aB���e�CAd���>���x�ױ����q����d�$C�]��n���e2�Gm����sN?Q��'?�hL��Y�ג��	|k�L����y �߼����{p]��j�D*UQ�5������U�f[.�&�N�u�AV0q��{�cO$9[&X�!I�ܐ�C2m�J:��b�Ů�{(Ql_0�E$���'���b���g��[������F��Z��Sw��o|-vL��hf^Z1�ҁiD{Nl98��}�VpϾܶ� �ݻ��sm�urh����st�ɖ��7�n�I��Uߩ<�0��8�j.��x�2I�V��&zݶ��� �2��6i�͋:�aLl���u4�R0]@��r���̏rUMR`���j;^O(.WS�Z��6�[�QҸ��$Y�<z$ �OC�a�W�}maV�Y3S�6���%���)���tk�����F�� �G�7n���ѡn�Q#�+jp�Oe�%*&1����^[Aku�n-�o��?�L���`��Ɨ��&�ήa�٘���*N;e'���/�eO;W�Cj���Q\�C菌����9k��:����w�纔�o����g���YPo &�,KK��}���}��Z������r,�5&ШObӦ�Xg�q�+WQ��ɞ&�<��ܐꮕ�^�n�~������Ѡ���<�z֥8����c�4SX\Z�]������̡�ic�t��K/ů��ը�b��>&0���%����ޕ �\��3����@�6K����C�,�ml{L����~�-?��?�s�U"����*��dP*W�\oa~n����B�_N�e����qʕ�d��Ix��K�T��7�f��}UE�:�<rꍚUن},/�᡽�`~� �{�1x����N;�:�Xl�ܤg7���n���⵸��=;(���_|�����0�7�o��p�wj�����$��[_���XR�AE��ȧ��(�A_|!����3Oڡ;�59������5_�	��V��he����'�n�gD�\{�X�*2�*X�#�S@g�p��E�LI)�	�y����Ɂ��{���*ұ�6�W������0o��d�R�D�K�FՉ	�/ȩM3�<`9kV��Q�X]Gsn9:��6j�l�D��D���^����w���2A#{LW����~�r���vV"9.f,Ɣ��6�p�)��F��q1�e��ς�eX��jT�SJU��hT����`�?���x�(��3/���e�>��yȄ�#0%(�L`,-4٭F��䕴���$?]�@�g�$+ٱF[�����m�T��J��"��D&N�:�R��`�w��/x� Y�����Q��L�}V%���[��n�H����)-�9��J��`53R�b�k$����\>Ӫ��,�`�ma.;    IDAT�%*��.Xs��g�>�[�#{<���E������.��M��~�2���$�Ćq>��6G�߇0��`bD0���^s C@��YsG'+#����x�y�H�{���Р�<�lZ��FBe�)�L��N��p���3F��������
�Zw�4f�\�#W���4����y�\=&o�ݦ�3)K���������ֺ�V��S,��*��I���&s"槯�of��`L�L��0�I*���P��]6/�$=�aޔR�0�S"�u5�b�D�+���}H�?K�[!F�D�i����5y�׉1X����刊$)֢�E_�����=�4��0�5�A���j��g<�Ѹ���p�'�QGm���EU25>�&}�^�ܦڍ���������=ܱg�^��k4H����6��\�r*��ϧN�m���;E�F�cW��ƻ�!8<�z{�?����% j�3V$`�1/\IqS�2�w��>��L���C)*��.�CS6>�����_�����1$����~����k�\3�+�YX��+�}�nߵ��zXZb�������%A�]2��*��dZĖ%So�6��ڝ
R���#T8���ּg��.2��VPۺ9�m��뻔��E�1�'똬T5%`en��Iq%�g_o��\��؊��)Imʇ�&j��议c���y��(֪��\�I���(NN���g����Zw�-qv�p.]y��8aۏ0?��A� ��w�����iw\�q1L�������G~ �4�9k�����)��M/�%g�@��97�:�?x�_���ݎ6��u��zSS%������R%���wx��?�o\� ��I��Py�En�Ba���������q�cL��_���_����D�?F��U�p��B����W�(�%���6�ШO	@��J�S�k� e"� C�i�P2'2&�Z&��nc~v�+ �^��(�I
L�H�3��rk����E4�y�꯼
o{�/�y�EzW����'���~�͏�Ec��n��I���E3�H�:.�K�;�^�a�q��~�7^��<�dT�����Ự��z�V���n��c�w:n�0�.UP��%�"@mLnF�F4(��`�24Ô��@z}�;�vZX_]¸�kj��\°��A���[��m�VLML�^m�5�}<x`�?��ᢇF�������o�YLM�m�:�� ���W�;߿C��x�O㪷�[8Ĕk�?���ǻ��k��6=�G���S���N\p։��,�����?y>��/�Tߡ�_hT�����\���^���s=��) ���j<���>���fJ>�����p�L+��7�pc䆞d<�p�8��r�8^�V#qO�yOȖ
�N�Q�hh0e�R픉�WL� ��Dsv�N�\^?[v�T2^4޿ă�w��Ȉth��K��$SV�0��F�ѤL#-\^��ZN�i�����K
�2>rŢ��qCڤ�ǔ�D�?�v��c�J�8���F�L	J��.�z��}�!S`��Ì]�P0�փJ��*sA��/dZJc<q
��Ʀ��4�bf]B(��7�1�u0 ���0�H�^�ԓ��|<���$�tgC2���>I�]:�|v7@���p���P=��^dz=���?���*6aVR���l{�@K�p�c�%E���tZ<1	����۸��� #�N�D�͈�\&$yћ�E;�|{H�}qьvB"M޸�Z���ͦ&�J��nͥ94�g��
���:�8����q�9���G�5w�3'ߒ�2�O���r�gA�]��{µ�� 7޲�����1��d��\��<l#�qi�X����8$��
��G�y�^4���`������C���@>������%��`�8���nY��]-�L1�v0�F�
_d�A�_�,-˩z<H�?�&����3eۣz�xhF�'�Ӯw#Ȳk�b�qi�Rb"��T�S�>N��
uQ@�ש0�j ��g#����D�:��R�Κr	��`gh	=ԋ#�z�N\z��q��ǱGLc��Y.��r�ҼF��.��d���k������Mȕ�P"@����_>����UL��bEgch��X��Ȑ�ț�{z��D�$���5x���pF3)Jm���+�$2�8��x]3�S#�4���ޔ
J��(���p���u���W?����2����`�q�������*�B�f�װ��:��=��n{ 3�=,7�h�1s²��$����
(o�D�Qǰh��$N<�ڊ�)01��Q����:������hlߊ��$����RS��r�%c:Y�D�"�E)/{D�F�S���Q)I�&�"�H�����5�-,bС�Հi���~Lm�_�Zˡ͟W_�Te#�Q��V]���oՏ���Q�1u`:۫�3*`D\zf�΋���(�t�l�a�]�i�L�o|1�t�V��c��ǧ?�u��?�����mYpo;r+N>�X���^��N=Vs#	L�_���O���߇�-���s�t�ȏ;�Gm"0}���8%�C�կ]����gqh~=J?���l�X�S�ʫ gW*Xm��:@gP@�ʦWS��ਚ�]�zh��-�J�
}�]��C�*6l�?G����y��I[	��m݌F��W��%x�3/V�H������#�|�Y$�%�d������zeeWO�<M�	NQ�CAR�~_R�
�)����^%ƴ��'�y8���]�A�t˝�#�����"�CP�
�^3��Eɬt?K�rU��eT'��J�_��UUD�N%>V릴��m� )���w�1Y� �1굲�+��&��J����յ5��4�������^s�f��K&#d�ox��߽�n`�ų�q��w������&߼�|��>�]w�����6^��+�y�c�G�X&0�ĭ�����v�9�1�m�ƜՃ�ɑ&֣�=Ҟ{X�2�q�;n	U��D�`U��W�U-��0�s����,Jx�Q�ꬠ�;�H|���ILGd'�(O4L��k)K6d!B����2����1�,���d[�O�O$�<�c�
3�Ęķ{��6[Θ�ĸ6�mƸV0�ʔ��̌F��N��pyX\A�
�6�Xb"w�X��q�t����n��zD���H���K�Yj�����@ט��UdSo����0*I3f"4_���Ak �$I�T�����HD���Ʉ��X9>9�u�f�g*E��1�"*#��� �kz�=<��75�hz�Yp�C,X?C�>z$aI�	�%?v���#�������Q�Γ�0p�^S������싕��*�oÄ�.)�Ee�`J�FH��k��W4ƨ�p�MmW7�&)�MF8�u]�ⅯX3��B��)�����N�y2죻����9[�v�u2��N;
�~�Oᒟ:�UA�D��L&nx�^w�v��F��u?�7�}3��=$��q��
F�eN�*����J�5�Ux�qͻ���Y�`;���ߩyO���B��� _�s{�W�.�a6�b�%J�d��:��)��r��5Yd;9#��G6e��B1଺=W?�o-Ύ`g�O��ZHI��}tI��|�$�4[���VH@����ƽ�K�kU�sK��^�=�#5�3��G�<d@�!�}��}�#�t%��W�^�Q;wl�E睎g<�B�{�	8jsQ���u�V]c��Pk�^96�NF�������×�~����0?�q���畊ZT�ț��RL��Wm��o���5�_���{�8��nU���~"�������V�lǣ5��]�E_r��Ҙ@�	�P�};C�5=T
=���㏨������\�t�r���,0�"��Az~��#�<���έb����}7�r/��u����<�x�cμ2b���F1�G�L���K�2��CZ'�`J)/�]S�S*9)�%0-M�R^�c�)1�T���J9aL-��36]�l4_��|��s/�P�Dl7ݨi\�'�1��d������MdPo�T)��T��s��9�ϔ>4\%0���%�%0��R� ��`:׫��9_��v� �����l��b����������wbBǬ����~��-���*��<���ގ��O� ���G|���v=��v�$)6s}i�wn��W��>q�I�7`i��<�u>��X9�ԥS�u��I��w`��o_�mw?$�?j�s���c���и	��X>V㆝%��s^}��8��M�̕�Z=̐H@�rL�b�4Ƙd2]�`˖&و\�E�����󧿁V���eF9���N��sY�o&����e�]�;�X����Z���`	o��W���8uap�1�#�}{�c�ЂzK%�d
�M�A�^�V�7��q*h��]��wn�3�]��8P�.�I'232�aO�>?X��F�]r�:�Qزe%f>r7�����E�C�z�'��Ul�4��[7�Z���iRއFx��7�~/h�}��G�C�{8.#!�����"���}�;�l�T�f�d�nՋ�]W���V�[��&0U�����m	qVD�RIOF�P�=����нV2��E��Dmf�x?PM��	��C*��P�vP��ٱDɤ5�e�:l}�2�*5�1%��\��;��~t�� �j�=��A��g���Ǝ���y1�>��@����9�,칠y�zK�S|� ���1�m�w;ck��=2�56㯬KL}�O&20fG�b8���b('䳦5�@�5�2^��2@�9s
�*�8+�T6}U�j�5cB�U���d;���gNC"ok$�i����c� �jlb�p���Q&�䄋��f��E8ы��Ò�C��sE�3ٟ�
�QG�n��x�, 	��$�^F*XUO��d(-☔��9#	��{A0�AJ����G����5cB┼�oL
��v��b-����8@J�i���ѥE��a�1Z̀�0{,��o��wY|�)�`�
{�z]4�簶p��9l�.�sN��.>���8� ��ȸސ�9b����{��;7ލo�x7n�k/�����^��-��L�X�9��%?�`k�t��p��Ix0j6�?��%�~Mzf�=R�f����C��c��8pS��0�R��yg%iFp��$������
KI&6".�u�,��o��б�U���9X`�m�ލ9E����~Դ �ĦÀi�e\]��T�pn�s9��ŽHc�EعJ�)OT��J*,�$+7��5�u��뚫;�#?�J�~��*�t����	��	g�����Q	QK�-����z.I1�nhyǮu|���_���_���@�>�b}�%�,ԳĔ1<Y��}�W-�>=�+,��V%a�Sd����:�{�����Ԟm�бж��4b��d���_e������032��;������$��p�Q5\q�E�򹗀���%��V��M�=3��O���/��|~��Cs�x��*�g�ߴζ��Σ7�����-M$�R`�c^8/be<c�R�!���h�
Z���ښӡ�)�ec�V͍g�*����Z�
���|�=�s��Hc�L���$cLy�&���բ)`Z(��bR�g�;#V��6`�|��kQ�Sj�>��S���V�x�	�x��c����_C{dͼd����(7��r�L�dpqU���-�>�x�9x�K��c' �����8�<�$M�b��'�r���k�ױ��\���+6U��k8fK�����N������=O,|��$�$��d�<�w~x���O���U�d���f���
e#�RAׁ�~�OÛ~�2L�}�_?�l6�ʲ&��o���'k������k�E{XALY ]�ˉ4&~V��H����oH��|��XG��J� �~Gl�9+`zų�D��Z.��^��k�Yf?��O=O�Vɮ�~~�?������X�1�א��:�r)4�S��Fy�qg�\p2~��_�mS@��ۦHx"a���~N�u��A��/v*(�~h��\��`�^�{-U����~�_�I�9��;l��n�<a�	n[9໻����w�s��\��b��>�>�	6���CN<RH=<q��=�fz����_U��&O�*I�ٌ6k�>��fGf$�^n��	�#3\� 7ʍR��Y6Y��2�V%�l�q8*ydL��-��Ρ���孶i��QhT��2�@ɞv�xKt�cJ`J�8&��H
�n�1w)/f��\.�@+X�Fh�L�����*���Ι���3��U�K5έ�LD� kb�\X� �`d&Hݾ�<�yi& &� @�-.Y����񐓞D�Q�򵭤ğ�>��&Z���������$=��:"f�WR�0��-}l�L2�d�_7�lĒ8��5�t�?|߸�#c($�(;&�k�Ihսs�C��f�r7�q�=�� �Dt��F�ėf9rW�HiU���s�~�GN��D>,9��xO��Θp1Id�/�m�pa0��fc���Fo�2evFz�Ԙ+9�5�����~s���Y���oË��\��q��>3����?�|]r��QP����}3���wo�u7��]��`�5�(_�gg��̈(�(8�N�.��}vW��<��
.��l���>�b �
jZ3��YI��ȼ�v���g��Ɠ��yl��&���~�9j#�T���s+F.�����,Hq�>����E�1�(��)F�z?$I�E(z�}abV����<��
ifB��ʅ�U��a�k��)^�@�1��~b��؝�.��%JMf?? �'C=�6Z��ܰ�ܨ�2z8bSg=�Qx���{,6���s?#�{�ؔE�ܘo�,��^w>�ɯ����#��bc��[Plp��H���M�C��%,�+�d�O�l���Q}��$�n<�x��ag6_��$�I"��%����b��7a�=װ�d@Ts�]����vL+�.r�y�|��|�O��<잲��Z����p����?��f�V����g�߸�6��ʡ;*a�3�%�
�$6r�cZ��2�.�!�`��Hχ�T<ϡ1��w��Ƙ
cQ�K��RA}ۖ�S�xIQ�i��9�,�0����*��fSJ�Y,6�=�XD{q-Ό���,r(֫(O�O��V�z޶��{�\T�E��f~�Ge�A�3��9���^�L�p���|�&�1y� QZSHZ5ƂT�+9+S�S3n���!�r�I��W>GNA]�G7A�X��d�����x��>�]��Q(O�?����`���q�\�+m���7�S�%v�O�K5��I]�`Ԉ�1�.d
X�����G��\y�Q�RE��� ?��(�9(a��:�׼��x��]*�]��0\ؙ��"�(^�f �4�ܥ"�;�򟾃O~�z��5tXr�Q&˞�H��@�a����_I<�������{
��|��!��yOƛ��tZ6	��{z����s>?��)�M�Y~��{��V{\C5U�X=�1r��H`�ޥ�`Ϲ�\��_��I��<3|ñi�`�b�*���1�}x����~�n��*�t�����]�'�y��m���j�����3}|�_��oܴ�<���̠�-��$��0/�RL��I
Bz�g���;���S!Oll�g]��� K,�$�ɊY�ǯ,��θ��o �q����SSvU�O4��JPmF�wf�)/��������6_D}�&ԶO��Ǌ�̅��E�@gb�;0%c�T�9�|�dk�ʋZEn��1�j��4:�L'�%�W`j��|��W��@�Șr�֫��E�JC��( V�	Lc&b��<+&t���L���9`���a& ���sU_nȭS3���l5\E�p2���q�@o{~��UH���1%��F�aJ#����ǫ$�L�fMϡl�����f��,���>g����3K��>)���5�f�B�e�	(IX� �Q0V�IY� ����$yl㬉�LY��8���Hm=�������1~�+��s��=��,SF�g�eI�]��{y�|�MM��9�2)�Ԫ�����PC����?�qx��.�IǗ������ǋ���c�Wh� ��y�|��p�{1�:@/�P�CT��<ڃ�dZL״&�<�E���Z%� �:
�0����za��S����'�#s��6E    IDAT���:��v�`bDaAI)�Ы����K_��2��b��������}�g��]�L�{)߳����P�dv_���J��N�\?hm�l}��f�@�~�8sByNr>�C�9�зqi|QW�xۈ���b�b���CS5��z�u�5� ��&=�Ml��p��'���=�~"��VB�F�II�a$�b� ��b��y����?~��m��S(56c�6�R9�D�m�TЊ������9k ӈmRx���<�������,I���aJ��p���/���,|�����S����mT��6�S5��<���9OB��'�t��2̮c�K��{�Сׇh��`2i-	Foq��S��j*|�7�35��1�G�cJ`:l����N���1r�*�[7�D��42W��T4�
y�����70�⫕ה}\LQ��\�S�t�^c�]^E���mWly�1��Q S�>�,Q���+�u-SՕ�����]�'n�{����`:����P���9֘1��J8��P����Mp��)��_;�M��}�9x�S���=[74B���@F	��:p���_>�%�z���	5�TG�e~�6
bL[(��񮷿ϼ�1j����oyJxG:��Ԝ�iG��H.��u�o��[��g�E�2�>g�0�.Q�˚�4�=]��9<��q�o�R�3�����׷�)���/���}�¥��>����+Ma06�h����s��f~XJ�N�/�1Ht?���s�Q���}=���iɩ��h��s���V	�C@�c����/�5�I�:�ݵ�zL�>���E9���%<��3��7� ���P��
_=�^J9g:�gjR� �wό��?� v�[Pok}	Ӎ.��x�eO�Y���[9�Ğ�2+�,0�w8n���~�|�[�b�O�2�c
r(��W�'���'R�@�m{{�-���q���Iz�e�}�9��۳�Ä�!=�oT��%}~���>卉��r.�q�����c:`��QSO��b#i֬TK�J4L��g����y��]�&��)Զ3`�t���(���(�80�1]_W��}0=bK
Li�� ����0ͥ�wH�Tݕ7�)T���Q��r�W��S�c8�ڌ1u�Lϟ̗Ɇ�prt=�@C�n�nW���X�`��5�4��ڌ����$av� �55Iپ(L���_9㉨^��i6yΎȬ��:2}m��G���M���ٗ�_����ӓ�0����`⻂)s���~��"�G��c��{Te7�]���:���?��?���I풎��B��A��q8�0Mj]�C�,0u����iY��2դ�dף��糏��h��iɄw���u�1n/���5�����eO{w�����6��#�W'9���"p�\������o�J�ʅ"
�I�����,2��	չ��� ���r\�)�8�|	�6��ʨH⺢`a�|+Tس6���v,�� ]0v�d�ņu��/5f�5���9a^[��9ց���>�xf�^��K��5sdh�*���2��;F|��j�]���J���|.o�%@ӎ�4���L��yc�}����� :����p)a��dךM�d����`/uZMma��g~�Ri�X�^d�g9#�Ӓ�硎�����T/₳O�ӟ�8�w�I8�*&�(+2��>��'`J=ko��_��v|��{p�bv}�|}+P�¨P˦�,��B�Z-̗"�u(�b?���b��P�<���bj;����n�i/�eY�dI�.@1�^1������*�c<蠔� ?X0}�3/�˟�d�'�1uC�LO��ΐ�2���b+�4���jK�+���_ĭw<�}3�_��ϡ7�i\�)qŀ��d�X��R�2�͠19o�9BE�ޑ0��v��ut�m���*�[��R�h�����ͼ��W� �\����%t�0c�}��]ǘx���g�8���a�V1W��U�VVd�V�|Q��8Q0r�r�5���7�ޡg�Mf�i�ߔ�х'm�{�J`J���1)�zL��s}�rL��'�f8���M�cG�8t{�]E~���B���	G��d��j��R�UP�������a�K�s���{p�@�������kj'��m��i��
.8}'�|�O�����e�B��a����}]�[��cUw���_}��r�r����0�v��IFCJ��t`}
���-ox�;���(&z��޸� +�O�b����� ��<����Wpǽ��k(��]�i�����D��W��0H���hX��Җ �A�q��.~�/�嗞�ֺ�x�9٬��2͙� u3�G?�}|�s�DUI�dh�~�xQgF�*��<X���(��o\��@�|� � ?0=���0��h���U��?�',�ƚ�ʙP������،�wnǱGo��D��%'��`i��;�y{ZBkH�L}1��x���-|����;�+�&�7�T�C�V�^�1�1�e���!��f���^_���4"��U��>m�	k�!�� �8�yE�Of����"Ɣ�$>��.%f���c���L�(�29���I���c�̌8����F�=����5�ф�o}�1������T��6Z����JG��u1�`M{v�向rM1���U�*��2�e�&� ��&;o#W<ySRD�+�<Y��%6��sv(s����4,��03L� ��"�(v��/}pي���� ˰��#�1�Ypj��~&a@�&�	�&��3�8>2F�6�����(p��C�2b�$�q�L�dA<v
L��}q�Jh��;����>��Y�/Йd.���Ȥ���{�L���Ia�^��~"�s;$����cU��;��O���î}��u����?w^�F�sJn�*�v�^:�Ҩ�#��蜓�~<{��vrաz�L{!��Nԋ`i���{q�����]����F���
�4/*����034
%HV:�y+2Pb�`9�����=���X�5a�����1��4�Y���V��e�enj���H��1ؖ�>0��{��s�E%����������>Bį)
�!�L>��H��#fـi��T�M`��-Oʬm��Š�VN����7��p����@���$��������F����T��t�|�V(b�U|<ɜ���3+�
��y��ۙh�D��A�n��*0l�8�b�2�	Gm�E睆�>�b�,��9�2cj\S$1�s��Z�zP�{�^|���������)t�O�Ẓ³��@������`&ͅ�U��K�LA%��
͡�Ko�⥳ڇ3Ժ߉�WRE���]�K|2n~$,@��G~ؔ�����W��RS���/S�5�Lg)�]�=,�����k�]��g�/`ȅZ c��8���P��jU�����on�hy�������w:m����ʫظ��d]*�,0eN�u����eS�aХ��Ձ)�`L����1�������ʪ���
r�-N�1*�@R�Ͻ�v0�����2���7��w0@���zoE�響�x��\�xݘ�jl����~��C�c:O`�+c�7)��$߀ֿdM��V�TcK̹���v{�q�+Pm��F�Ӓ�^���29V�P��%���Ѐڪ�����s�~���Y����bs��#�OcǶMغi
�J	�j�rI,��l��lH=?b9؛P��zs�k�g�,n�{�!�t���q��<6g�Xq�n��@��S��:��y6O7�i���<je��.�YJ���W,����`��þ�y|��[p׽3�*F���@�?�0��b��И�߂��D�^��8�f��~6���_���-<������-S��l�~_���kt96y48�3spfi�O��1ڝ:����| {,aT �������!Y��ޢ>W_����c<��pޙ'���0ըp���������	�]�%��}\���p͗�ð��h�w�D���A�#c��d�|��X
�')U�3@��bu��$�3^\	`'�A���$ �ޙ-�s��ȵ,����驁�񝑐yT�R��%{`���p�a��p`�Z�ot�KX*w��}̱�8������S��Y�\��&�]������VC2��T�L"W%��}0��8�Q�Tt{�,��jp|��BsL��pT�u��.%����õu�QОݒ�0�
#"e���,P(-�Xe\�얯o}�2r ��>�5���1�v݁zN�]J�Ӟ��d��!;�Dْ2�T�hx��QX������1�)V�VS� #;�2zH�ր��Q��R&�1\I��tc�z�\ؓr�������T�i�'���4ȾY⊛���K��%��2�O2^�!�ˀ�G��?YV�&Ŵ��0�6�>���i!`�������9����:�J��+(����j��3���ݥ�<ͻ�M�P����5<��q�ǂ���l�����p��`,����j���E|���p�M�03�ĸ8�V(�j������d�v��Yh)FlZ�s�.o���_0a��H&�;��qc��:T��9�G�#U(�gU�&� �r_e�ڦN1�.a���z����F����W�����'�k¼g���e���?2�'����B�>��:W�Lu�2�!�a���f7π�̫���{&�ޯ1+�7�.�)��2�/����xq���i����#��LTU��Y+i��U2n�����v[ȍ���˞�
�8�i<�����˟��5�)�HR�s�"��� 6��7�GZ���}3�ׯ���wp�=s�7v`\�8e�f�2��ט�ډB��u���jZ �i1
��8i��Yl�$ٳ$eN3y�
��yM��p1�C�>ƽ����,�9O=�{ٳ�S��a�����?S~��gKu��r�ְof�>��[�z��cn��V��yzF�����R���l�¨Z����֙���X�SD�1��\��AkuU=��A_����9�ک�c�^�G�����m�"s`��­lR^Iqe�H)p����ӥM�Y!�y���DU�iHg^�%�sLUl�x�3�]�S��*.8a�BR�ɘ��ρ��_`:�+o	C:�)�MB�&���2F���e���A��>J&�v�4��4evy��T��U:4΅��J+����0�[���7�d�
Ͱߑ5���zO�\dy�!�,Z6�'(��X�; gVP�N�Z��{��4*l�"r�Ǆ��@����oa�YƠ��2�S��ۨ�� �G�@�K�M��>�o��r}
��$ �!��ؖgѤ�%IZT��౱��n��g�-Ü�K%�:ml�4e�%0>o��:o�N:c�s�X�ܸTA�6�B�sD��+(T�����9�$�N�У�_��}������aG >�%/ެm�DF5�?�{�*Ͽ��V1����#_ߌr}2�BJ�<��m9�5�Lm~�H��$�yv�3(���?�3F�cn�&%2S���K��'"{(�6kzȧU���l�{2�\�3�ى�p`�rV��}l)�׈y��WL?#�jk�h�sV�m$�n�/�jf�PU�5�%st��t��6��*S(o� *%s���ƟS����z1^���,���Hk��t���[�ZY�T�b�ۥ�*��@�;&(�M�����%����Jz1o="�Z�m�i�f��^�#r���$���񢏁�
�v�D�nq�^/��L� ����l#��iˀ���f�T)�a���R"���8S��9+�JF���#����ٖ�7��g�]�ֿ9 U�&��X"��\����z�62'�E"dIz��0�J����ۗ�u�����c=���ƻg�H�2oL�q*��TiAƸʔ����0V?�?�:R��}�vئR{KГ]>&K��x��p����Bke�6Up�i���x<�t����\+�ً�����̭�X��7ܺ��]����q�|]m'<Ӄy�Q��{��_�;i죵7�(��$Y��O81�zm/�`�P�"24r��,�I���֟��C	H��[jb���.�T��X- 挽��Deî)[<�Y��Ӝ*mb�8%˛�my�<���q�zC��<@I��`�m�gv��lt@Y��*q�Lv��o�k�R2Ō��g�}-��˳��:s~���O�QN��H#��H��0����ԃ�6����nS�q)h�D��>}�+��Q����[��<�=��8�ILPH�B���K�f|��~*�@�ܽ��5��7���:�kq�%AL.�J��"%_̂���\�k�=�"�΅��~��D�3���K&�d|&	�j�:h�F�K�Q�M����~�zbL�E�����3���z�zLe*��I��'�����b̯c��e�o��:�}�XX�ӧ,֌�dIS9����S6�J���,�S��#�����\y9�4L�1-���S�1�7��#�ƴ�q1����[oc��* O��zY�C�f��W��ߗ�w�^C��w�=�ƘJiõY)�1ئ���x��|�r=�OL-Y��(�Vq�L��H`j�(dL�v�A���鐮��$W�l�\13?b���}�߱�M�d4.TJ%8G��� �kr
�[�<�T��LE�f�C�zʫ��T���Df�αj^'�����Z���
r����LN�Z+[�����#3ZR��"�9TA6*Ҥ�K�T	f�q�s�v�Kh��t=�8+h9���\@<���q,V����h�'�x�|Д��3q�9�ke���yo&�p�%jfN`�"�����{-YL�e�G�=/x3�h����H��gWA�`���9ѕ�>�de��z3-����}��M9�88�r�0�����9��ҟ֍>{�Xyd�ի|	��*�	}f�?c!7s��~�f�Z��9����]��.|�E=" �>_��$��#O��&;J��LN���Qm�fu]��h���U����e[�0�"Iߌ������h#�7?%$d&)��X��l.U�� �
��c�Pfu��FoeU��E��n��a��鼣,�}�XM,(�vW�4.f������9*`J�-{}X��kHʛG����H�Q�1�Pe�-�"`jN���q���/�%�NNH�K`J�4ƿ$�C+\��Ƈ�x�#��}�;]��mgl�I�dA�Βa�r�X�J�5��Jx�ӧ8�r�K �4��0Y�Cg$�i��V�C���		 �ϒF��Q4�Ղ��ԛ�@�@s�]J�=i`�^��8 �����I4���Q�gU|%��Ѣ��+	 �[�l�j}�ػiM�P�a��l��������5��5����1>[�R�h���)��~�gcx5�`�Y�cOމg<�\\r��8��"�,�{a�+�]ɳ�_8�q <03�W�u��i7���(��I��5t�W˳����@Hg�=�n*Y��횙�H�~&��2�+���s���ݟmJ�[��<q����@8$��&R�̜�`	�k(k��;�b~��ה��^��y��7�6��Za���v�Z�3
-w��'�$�F�
��&`��;^�@�G-���M��3r��}-���e.���\RXI�[���Lߙ�������n��������b�±�g�@3��>d�Zc\������{@w�tח1�5Q+p�c���O:O:�4<�1�1]so�`u��ydUo,P�~�!|�k7�[7އ������\��	s$P�h�M��w+�J=$7�k�օXc�=�0z���a�r�&l����9�o��Ρf K�;�����^�O_t
���/c�0`����������oڇ*���M�̯��}����9ܱ{F���}��p�}I^�m�(U&�TON6��WJ����2�c��1���6WV��u��X�iխ�d8ɱ1)�p`=������̬������L�1���^�1mK譲�t̀)���;�@O`��������#S����́����o}N���b6ӫ��,j�Z�*	e�.�G�`J4�/ׁ�}T����H��>�L}�#`d���J��h	�+�Gwa�����d?̃N�H���fe�mU?��]X���uhZ~6    IDAT�>)5��J(�hYo�^F�'$V�*���b�OڧB�\�i��F��{ۭu�V"��P��Wd^���;��K�**՚�7ʍeT! ����@R5��vd�nRLKZ7F+�����Ju�b�m��F 2@Ϳ�xA�;�#6F��I����l��c����H���Y�V�Q�������� �Ȟ+��}OU8JDؿ`U\a4�!�Y�U's%9V#i�S�؟�Ƈ����M��\�~�(=S�:���{�eS9���`����m>� �M�g��UMݶ>��3iUù$��e␈e���@���i섽F���� ������F��	�z�t���9�L2�E� -�ip�W�������?�N�wK����议��j���S{\O��,��� )����t�0��P���Ď�UK���T�z���t��ZZo�;��9a	0u6RUA�`���(�k!জ�<QG�="���i�hč��l�(�.�G��t�H�Kp�X���0�\����o�W?MJ��j/�%�?���u��ah��c�K�"��a�ޡ��,w�ؑ�ψ���d��ia%�#�"P%���Pf�.�������z�yI�A�_\�|��ߗ\h��M�!��>ds���<ςbڝt�.�a����S�^���F,�Z���<��q#U���K��Fa���}J��2B���s�N����*z�%L5��2��S.:/y�S��EL�ǍkЎ�8���>�U�;7ދ/}�Fܶ�V�yt�H���;ز@�<y����J̶����-X�x.ג�G��w����~ļ�gI������h�(U��X�.b��9��\���1v�,�X�����@J�2��E��b2�	���
�*jZ�dE'O���;���Ե"eS̶��f�~-���ѳ��9.�Y����q�%2P�j��
�N��n=C�HPrc����e���`a��3���B��Lg������/QUy�[�~+�GQ�
e��
Ubq��kB�P���`�Y��u�8v{�<�4��YO�'��D5�"��-�$��JN,8�|��~w���4��;d�8�^��׌�'_���e�� ��
�l��y��#Pʄ�tVr�������`_Oݯ#O�zt`Jƴ��"7X�έ\|��o��1=�&EΟ`�4�)����bLw�?�;�ŝ{bf������$4L�I���Y��S�	����21��(�򠔷Fl��`}em��Y��V�zL'��	���ոN�N���2��̏���Y����*�'V�S�*j�c*`��~�g>5YƴH�4�i�ә�?�;Y)�����'m�{~���50冡�������������c�"ࠛ����-�	0X��т�W�&�z���$��+�Ѥ~K���܌M�#� �X�ѰM]��
$dTիh�*d�6���yx)��� GF�q�E�r����D|Yҗ�Y�?��Ƥ��y��Z6�����9�Jp���`�$� �B�bK9)�'FYK�����a��2���bG(��R�:�ʘ�:�HH �a���v�d�p�+&�6��p�5��?@�]�9R�3/��_4�]�D�sg�{�$I��+����� ���b���Y�h����.��b�^�g�9�ݚ��P���~���H����x8���P��{�<�4�u#'��g�Yb�:��?lT��R*�L-I���Ȫ�`�Cw5̺�,E).�0�!�]�'��*QE_��r�IƲĂj����2�M���Ө�1e���$��%ܓ��r��/�(�YY��Q�ד��R��#L����U��0j+И{8�����:zK(�G���3�[p_c��	��XS�_�k�]�ɚ�M�'9�����%eڋ�������#�9�4٠*�R�#3J�r0-�Ӗ��'+��-֛Uĭ�L��d7w��>��@����R/6��|��^$y�dg���]O7�-��O*Y������C��˨zD*d�#����"az����`� �taN����}<���V�ݗ8�lK��F�4�#�$������L!ʊ6"(4�D ���bRV֛��ٿ(e��D��	�&�W�1�71�,c���Ӟx:^�����ӷa��m�Cj�_w�C9��ӥ~��|�?o�M���0�@�6����?���v�/��D��0��^����%����:�S@h秩|�<�}J�X��dq'V{�<��5qfM��Mf/�S4_3��	�zP�}�afB��Aފ�~*G�3�I�ґ$�7Xʔ1�n��P�������a�$�WN�L*�?�"Mܫ��i�۽*[����=L]�)%rc�x�y�}��$����ѧh��z����8)����H�S���'��Q���Ef^�'2>RK�K����Lz��T�]��w�ˈ1j�2�cuqV.����(tWpԦ2�}��g=g�r� *�����ޚ
'�èD�{��/~_��-��`����i�H��yxq�Z.e��m����"�lm����Z��������]�m1>��|�B_X�%�9��4�1�J�:9�u���15���܉����ǖ
Pqgc+���')�۝�%�����7l���Y����ݱ�W�̭���5�y�n�u �#o�����*=��@O��>g<�ع�	����z_��q�s�ݕw���(�A�#)-�N��� �$L���b�6m��� SJy�.���ۛ[zUW�����1���, 1�X�A3����L��������?��QUvuEt�#*����m��.\�a@F�B�ӛ��ݡc���9�Cu�;���޽���s��k��>Q���ŴmACG�Z���B���k�į9�D'�����HR^̬�Y]D�hsP"���r�)��0?�+��@`:_@�30����S����)�������2?r�jgu�%���ƯO!P����=����'V1�I��$��Ë��#���d!}�^�����J�W�3�i�x:���!`A�I�Ǳb4}�.1�
z�2H�yz&��m%"��\��#�'�xS����-��坥 ��N:!��wpV/��? �}(t�� �@tT#^��(`in���Y��?��d��d�F<���2Y��['A!�C8q\�i�Qo!�h��4L2&�p*#1�*!���HFD��
�e��x�M��C�;�s�>�{�K
�fN�5'���ɝ/����|p�
�]��q:�t�`O
����KT��S�E���2��'� +@~��a�$"s���(?������lA)��Ύ���`�z��� ���3&pt�̉Z�zc�Bʻd��]J��*w6���lR�{��i8o��#��t4����֙��1k$Kۼb�P��6�JP5'8���~�#�TS�nP�Ik�{��+N��U��y���g�&�`|���0ɓ�T g��P}���tp��D����{RaE����5��G�q$�IIN\�[F� �ź-+�N�� �W$?q�ٰK���W�&߀��:�G��F[�^-�q�S�e���Hy��� !�D H�x�"�J��3���^�
(*�l�
W�&; 5 �B��#�3�.���TLlt�k�����W����-�η�hW�6����KG9�ā)�.$Q�#��h�~����/�k�͚�6C?\�0�"�0,T?i}�|���̻�W����W1�$)�JC��k5���>D��h�ڵ�L��\P?�H$8q�3ˊ`2Zoz>��q��i��y	϶B�A��|��A$Y�>+_�A��O|0	�Xn�~���Qq��^�f8�4�T`���_1���D�%D�a�u^e�+r�E�ͣ�?�L�ec�Lqw�rpZ�AlK���] *�C?�J���R��qbx� |���z�y`:��&~����k:�����x�5�C�|�i�����{~�M���%���9�3$���Pev���?�y���m�X�icլ��t�ak�� �X�d�����.f��!�A#���'\
��;��C|��O?
3�M�JE��lzd6�h'{���Oٯ��_�]s�:��:8ͱ<�Μ_����t��\�Ϗ]��z
"[#���g;u<u��;w`w�I���g��������FUêFz�
�6��[�	b�e�k���s:C�Y��
S �]3���0b\���ݮ��٦J���x�v4u`0��ڳ�1�+/̼�����赭���ΜFy{L�zm[A����wwIv�\���ʊ�8.R^���i����^���s[L&֪�R90��`��p/e�����XL�5X1��ן���wf��5�0]�+V�E����R >�����
p��h.��a���}��.zx�2�ȩ=��qB�(�+�&��Z:dR��Ӂa��g��>���R��>{b�d������LԽ
�X:�â>�G�6�^	a��~q#��-6q0���Ï������R��OKy�����Fb�X��As�2���b��ȍ0����@ـ&�d%-���"ܢ��Tgy���%*����rq&��@r}��'�	P6�{/�v���$pq;i�Ʌ��Z���j}6���EG�[���	C<�21��Nk#�Oah�SP�T����)+��`#����<?$�>
�sf�����=TLu膳n�&��h��ِ?�ؗ��u�V�lR���X�d���]�'`:B�>�We�����3�cڲ�>7��DsF}_!V�@	�cG�.�Z��[�	m��i6%9k�~�B��e�S��B`fr]$�,��w��J��9���ت����P����s�Re�����@KQ	�3��ʩ>�rp��8�,���n"qKFZzY)�⸿GN\�+�P��{RT<�/��*���v��|��Bm�Sn��q;���,�xBIG k�#��'S�	�aw�gm��^�3���$YRb#��%"% ���@d�[*�a�� ���\Ad')�����*U0�S�<�?k+�����o�_x��u?z���$ۍ_I2������y��ҝߦ��#O�ZڶEs�9 M���$��s���-��ų� s��1`d�1Z�z�<(̱m��U��>�}$�i���u�&ɂD��d=!�D�d�/���ә��R��cI~��	 ���>̳����,��R���}�ן$�\r�`��7|H�q��x�s�W��cGE-�#W����{���%�~T��b���F���a�]t��<�q��EU�gcm0Z��_ݕS!ݽ��L?���q���SW�Ē6b�z�+�7}�h��0ut�c��s6;�h������-oy���g�lϻ���b�M*S�Y`�gv����{���۾��E/�9z���o�;�U(<WT��3ë��2!ޱ@�V|��ց�&�.�M�h;�s�
�����X�\��j���r�|h��E[o�����x����m�!9/3A/"E܎BC�R��������55�x���^~?:,WfO�ݷ��޳o���}��g�kzpg\̇�īR?S���k6ma����he��?���jߞ4ǴV�.r�����k\�l�\���Y��s. S���9j�H��
<�#�����N�Hŕ��{��pW^WI���FŴۖ���Ȏvwl2(l�@��Y}�'y�O)��W����ck�*���
�Xg6��d���rW�La~��;�������|�ր��� �{���b���i� G��eP��<'{
�0J����Gb��f3���q{�3�����?W�ܑ1�r��#�aQH�'�1�,1�<	c6�zM��y���Q�Z`)����+�d���t��q�	ƿ;��嗽QqX�����\W�UT�ԺiC,����3�B�U$�y�Zb����Kr�t�:�t�G�;LG�X��ڽ2�6Ѩ0��k{i�a�f?��q/8ܹ����Ö�{%H)�u������D�QC�~Ir��k{=��X'ma� 3��}�5-� 	��
 �i$����!�X!s��D�W�N)�]eS>ke`�~D��蟛ϭ�`;X�A�*k�Ć�\vҬ��_�r�F�HcfZ�OEs�̏���6E�q�Ŋ������a�h��g`
�׻�ѐ��Y�XAmѨ ��i�=���^yZM묭��G{��	���J���D��I*� �0Sr8�j8��fH�Ѣ ɘ�j�b ��^��n�u#|� ���N&=�ǔ� Iį�j5�W)��U-Ul�o@$=~my���%2�4w��k�Z\>��k�[��"�?���8��2oR�Ṕ�/S�RE�����T �[�R�b�}I$������ĞKyg|I���<'�ܗ~f���ƜK�v�BBy�H-6��-%Wr��������MF�V��է{��w��nyӍv�i��eF�J��n�qOs��}�w٭u�=�̾U���l��=ohq�+?�8�$I��*�F��^�-��r|��ڻ�EXNR�`T3��qT���4a�n��7�E�xE{E,[��ry��w��ӯ����}����8�ji��&k!-�y��_-�%�`���$���7ul&Ul��+��/>����S���k�3���2��$����ߟ���Eœ���]�˜sġ�FI���SU��=�F��WS�B�4��4K5�j@�80�XJ�ઉh(J�f<�MF6Yu�k��gm>ڱ�������A{�+��Ֆ�aϕD$��.�1e�lol���G��y��۾f��	��7��]�BHjLy hPU,`�(�U�oq�KX���;��?G%�k7�N�p����=BU���i���M�;֫�Vod���+�~�g����J��������/0-����"�jv46{�v�g��=i>�kO>s`�!T�-VT�w(W�<[������X���iq��
����&����S�4�)& ��׳Ωm��¤7p4�p=�l0[_�̏l<����)۰Ђ�jr��Ҹw�0�4��i�
�Zoתѐg�L���:}Q��/"Z8H8�D���Asl���:�]��lٿ��8.f��D��kO�?��O���k#��b�
x�"�i佞��}2�*��I���'>W*���O�r�$��tJl�K #�Kv,kTc���JVb��D�9@�b��Q0z��
9����x��4K�xޔe�>�C�IrSVS\��X�8!��K��Kp�!+`��P���,@�<�.���^���aw�:��ߣa���f���O�`�?�gi�h%u��:N�z�7����{�%/�X 	�j��p�̄�3*�.+�n��C�5)3Iy��Z��c��$�qgEV��b�U[�@?�#y�d��L$�d�3 �͌f�xKU�8�*C~��x��Q��R�?K��d(�������X OܗV���k�s��	������e�п�o����B�1=�i S4`F��SVџ
)/r�q�`�����m��[9uR��6��w��$����S ��a_=�3 ��H��ຠ�;
>�4�&UN�8��}�A��}�^BE�͢�����țcp�df3��֘�| ������J�B?���L����k� �s�N:�)q֓��]'�"�NF#i�)$�\�y���'�3!���x"ьʕ�x���i�GTq�t-��Y&�A@-��e�.3'l�9;����7Z�d�Imѓ-�λ^�(�|�T��]��?'�
5�̲$���C$�bj4��f�/0�kr`�������G��S���U��}���	%�����fO]0���O|�{�=�]�Ɗ� �`|��lb�>�ɫl�	"������?O.J�u:���jX �Q�)?�%�l�Y��!��E�^����:?�rv���8��1�#�}�-G�3���9�[��Ig�ΔR�.b�	���:`L�pA��s<z0S�5���L���S�&����������}���=���لG���������%u�RHɠ�_Pq�8�5�'�C	NS>��������>>s&{��p"�xfr��R�Jla*��jl6[�>�X�j�o��Z�ٻ~���w��^v�6ɢ��Vt�9�{�lh���M�����=|vh���9��8�"DP� m��|����R����r0�CDN��#�\;��⹅JE}f�̸_�7h�����&Э    IDAT��9be�Y߬ڵ�ơ���'�W>�.{�_l�(���Z��*�70�O�z,���Lth��p�����'��o?f�z�Y{����]�p��C�9���{b�����jX�䦵7׭���ظ���xYXf�f�J)oͦ�C;B�s<b^��J�VΜ"�
�]��}��O  �zS����۸?�E��#G����^[���)��]Hy[6*�)�6\׻]VLL���0��^��b S��Y>�X{6��h���B��TM�/��A~�BI�w>A`
�# ���K5�:
v�M�F�����v8�8�tt�FZ����XF��,'G��D��L��nӦ��cM�E?C0��HQrUn�\}*{*r �Z˓/��MzR-%x��OԾ"�C��Q1�\^X^UQM���KZ)�}��Fr�**.KI�u0X-��;���>F�G��WI<���u.��`��Qq
@W&��^q�~:�>*Qt� Ž���UY�9&�BԪ��l;�t.u�g� �VR�$��?��8PVҮ��X�a�ĵC�K'�7�v�=.���rc��GK�3�Ku�eh��2܎<*��.ĺn�����
[�"usJ��p�5Z���Y��o�v�ֶNZ��%P�~9� ��c,�H�G��=�5Z��ܴ�� �M/�6q`JY���1`C��Ӂ�)*�0?0�C�w���;�)	�+��* ǁ�H�
P�����g��2�B&{/� �c�qe�ɘ�g�>/T3��=s�ku��ɼH�bar䮹E"ǵ��%0�gi=�f�Ɨ����Ȯ���R58~P��8��lp��p$�E�c����8��h�H��=[���5Ii��4o�e9/_��?��)v�n*�����&�$��I �{P�{�Hڙ����>쉑aI��R&�b_�3c����Zc޷W��<{�[_co}�v��vs��jB��ka�?2��]���i_���vnb�ƊY�����>��o�R*�DD��r<�r�N���Z����x,L�T��DY��:�����7=O=�KG���?&�^��m��9R�,I�Q��Ɨ��� o"���N�i��GR�����4Ӻ��@���^N�\w!�*!�z��ęgg:?|(V�s"�$��D�@~�WRI�����Ahr�-�)��^$�=��$�( �2 )7_~ ��w��Z<4�z�p<kV����� G��:�+�e\)�+��h�Sj�T��C�����9�	��-�C·����l�~��W���6{��7ڙ��P��Lχ���t05���}���ߴ۾t�]8�\̞5Z+,@�����u�٧j�J��b�Q���F��*
���-H|M�Iq�#�X��U��!r@�F�}�d�9|vm�=�k�[�ޟ|�}�]o��.TP�~?8Z����������������ϑ�+�hR������q�w펻��h�綷?��n}�v S��$��&����l�L�V���)~����Y�V���1��ǔ�NF#zo�0)Ӟ*�x���X�Q�bf�+=[m�83~�w��z 18��@��bv�z]e~4���i��6mt ?�=��c�ƚ���j���5C��*��Ѯ���[�/~X`��O��c�[��Iۙ��h;b�\�N2.���A`��,6{�4gsG=aOO��*��u�,'�Z�W���WҸ%i�2Z�HTIS�^���!�މ]��NQP�%���|��.���0��}�R��J�Ti*eƩZ��"��R����8�{�f�?�%�g/ٿr����SJ��|A02gǤ7
��}E̈́!���H˰ �Ā��ĵ����!# ���Ͽ�ڨPFh�	Q���Ƹm�$6�z�V���4�ĝ��2��"\
���Q		��L$�~@��$��B&���=�5 "�'���I
;�"�	���-)�>�ԛ6��$*p��S-�-Y��=] �&¤���]�qn/����6/�i�;��?��Ĥ1��po���[�� ������k��f����ɶk���b:� `
�����G�3�����ݝ�e�pyn� N��aN��A&��E!�םg����RM����`����$�� e~Z���zOk<mV�P�us4m�̈�c��d��Z�"�=�e�֦?�2"GES[L�:bD _�v?YZ��ڒ٨��E7�q�$�i�boĳ��p�ҵ����W�A��ފ�a��_�Z�6��u�Ջ���;S\��5@2G���Ϣ$Z<�tH�s���K>���y;����6���y����{�KN��:9�F��Zi�=�#3{j���_z��������v�Z`\��u�3'Ʈ����������ƚd��Bv��7��FZo��+�|��s����2��)��OA���U�7-�-��x��o��t"��|�&�;��Et��؄��l^��&�n����_�%�H궸��wM��館����I2�؜��5����?@
',xU5�P��gG�S)��Ez��ܸSuU�#�����I&��^�v��{�T`���J0}��K��2\�s6v���ϑ���M|���I�x{�E^�@�T�2����pF]�b:�&n�|b���lڷ��m���M7��~�g�l���J�a|�ZV�)KF��Fe�3{�=�����_����۬�i�Y�V�69/� R���-�Ag&cX�<�� 阚*ڀ�
�����+�q�D����f6��[}�g�o��ꅗ�����K�ݲ��g|^I���Jˑ������lz�I�Y�2x����_���殇��wm�`a�ڏb4��K�`��g8��k�lek�Zu5a���h���܄)�-1�Y���H�x^��R�ۣ��}4��_'��!E�R^ Ӫ?�)-�G=���@I1��Ї>���n+`��j4�>i�D<*� ����@U�b��]i���Ω��*�������?0��zL�����_�ѧ��l���2��8��ӭ������gk��*��Z����h��D,� �@ɱ���}anF@��_���UT�ү�$ F��q�0�0��Q�z��X�G�U�>��6d���*�<02{�c�`�Z� �����Yk)siF�kVy��%������k�����V��L�&S�<�D �A6F�Ę�?��[u���ϛW��*�T$���ٱ��8��`�g���� �:}B��Aɓm����d �ʸ׾��:9����.����ʓ��M����W�3�3I��饘��L\(�*��1��I��^���	����2��.(!OAŔ���Ť{r��6�fM���Ć��vxp�Dx}����Oؼ�>JVL]��3��i݁)�fՔ�twc�VO���\ysJy	L�q,0���C���,�H���%�j5����$�z�iʗ@��ߐ�tZV��L%knh�%�p��z@�n|uv�i�����
l�i+$c�'8�1�>�Á$fq�'��dN]��� 3�{Od�f"Yk��40���l$2ULl��U'�3�~�K�l	D���y�ǖ�T�Mer�Z ��:���xI��r��?��|�R?r��f��đE�W��.��TF�V�������HXRYB#U�c��d\���3v�ɶ��]o�w��:{�5Mk��#�X~�%M;f���}{������w�8��#�um:oX�.�3�7�%�yK��}/s��x��2�	�
@�����3L����qv�%��ɒ�NZ+ sb���E�G�F��Kq��F��ڪZ�~.G��5������ܐ/~��g��/����z���r� V�=�Z4�@X�0z��ҽ�#�ǿ+� 0���c}=Z4�?~�x՞ͦxiE����}�9�{�5�Q1�<�r�͋���qP��$�l^_)�^<v�ҕ�Mp)�gI\g .�G��X/o�a���L��.^
�0@SE]*�{�5n��t��@����8��^�a?�?f~�;�,|�'
?��J�~�T:���}hd�ė����묝�j޴z�k�����S��…|wY5s�O�0����u�^��pଁ�ނ�c_�;�]2�Yud���6:c�j�o���ч~�6;����{&���q�������hT�B�] ��72���������������f��$�5�� �]1O���V�V�Nr:��Nc�)<D�a�t���ʉ;#��b���^��ڪu��	9���D��*33`Z�Ll��G`
�*�S$��Ho�5h�Ċ���Nۺ͆��v�#`�x^��b�X�ѕ�[��~l�9�|�%>z�1����^t�~�|؞�fX�ųN�� ��7ڿ�����hW�FG=B�v9��\����;/ �!ɐ���Ldz���cajQ�
�@q�ܴF��+�RJ�zU3��8��䇒�}�v�t-�49���+
����UPo�A�~^����m[>,"�/�� ���=f
�
eV�F�~:An��H@�a_ ���z
�w'S��/�dY~�|�9>w�,���]|��o%'?ы�9_4)�g��5�hʎ����%.\�R/O_�ayS�n��@���L��NmI�[��|���GB¯��sW�W%�q0'i[JÝ� [�D$=�[ޫ�I
0a%�.k
��l�t�7��0p9Ƨ����J~�`���F��v��Ǽz�u�7�V[,`J����ӣ݋쫨���)�V�0�	�د:5K0�+����g�[s:�^��+��*��ۭ����%������� �4 ��P�m�N�RH���I��A�=�x(F��������L��NY-�LŰu�Ke��7Tb���p��:bb����,�	e0���Ӊ=U�Ty ���Wσ�O{��f��$r�cD�H\�{��$�߈�^�*MacJ��B� �Q�
��UF�XC�8?gޑ$i)�a�~� C�Ns/�+�9�H��ϰnI2Φ6�_�V��Zkh��������nz�i[�Y.��dwAp���.����}��w��~���/l���v��(�/��ׇ��Q�Vj�>Ǒ�jѾI{�[_<�R�JYp^K>��x�A.@�T����X����`�20�͕�Rʛ+�`����q��^��*!?�4� c{ ��S��[��+��7 �]M�̂2���r�.|��^c�޲�޳�l\OL��8��R�,z�� ��[�F���L�`��rΥx�9_�yE�r�g�sy,I�/��XK&�~V�A�\�g'���zq�į�#������כ�6bZ�W�qdNV�\��Cʪ>b\:1�7I�'6h��tt`V���]g���7��"V��gNp��г�٧�#�O}�!�?���v�w/Xڵz��5:k�[]�4��_Q�ĵ��w��STs�I���gM
%��ySv��w�9�M� ����zge��1�Zeu[m�o���]�մ���%{�W�:H��w���ㅑb����k�4=}M�7�F��RpV;�����sC���kw~�1�Σl��	����P�����Y>�Lʲ:g��[-[;y��� ���K(�� �;p�1>]��`h��C��^�[5VW�{���z�4��h\����60� ���؆�����F��Վ�10S�VgX]荗��t�մ������h�Rޚ\yW5.f�ʰ+�D.�]��)Hyg��TSJy_�m������|�;��z�]��l8mp����63>���n<�d>��i1�!����1#��w)������+ gT�tH�[b�Se��|��s +#'m*�M�g@�+-��J�W3��ܥ^���1�)����p:��U��m�,`]@�7����U����k�p�;�x�4U��x�LJ���Ro�˓1�JEu �T���R%<���G"y�T�s��z%�_;�1���� �	���R�;mVx��.��Z=�WVU"�y�hb(�9��A�A����"(5�㚎=_׹TPTf#-Iu����
�6�L8V�pA��	�{UZ�I
*��27*��]�:MkaX�%�T�yS�fu��`�wd��C�*+'6
`��]S9�Ơbڨf���\�t�ѱ����}��+m��~n�3ո(�
x�]yG�?{��өuMks�S�����tR� ���'�A")�@�	s�| �-�]������H��[�	On��Pq�Z��_��Ě��� �<V�qpb*��r�i����p�|+%�K��1F�(�H��>��ob���x1����+���t��x}��C�Lɯ%��%�ګ0k?�����L�Rr#�"�r��Jc9ъx��ɻ�R���#��Z�Q]�Θx_�?���s��VJ��s0�2���)�®��]{����]o_}F���ĵ�8�&'nn��������3w|�|z��5{�6GJXǹ�$�����'�W����U�)}�}�u�T�+9��t�<N:`܉`��4�q�@J#��z�����8@j�ƞ3��I�����R�BBu����% ��A�1n@�� ΋83�H3(_�a��x�owr��)�óI��IO�Y�k�؎�^Y��Dh��XI`ϕ5-�w�?�������R��q���L��I������	�,*�z�!�#�)ymq=!	O�G����>�bz�p�����}y<_8�J����1�G#�MT�QA۴�hph�jdU׮����^�
{�-?n�~�e,dQ޻���rF��:����ٝ������_����vu�l\f��ID�.P@(@D�E�H���Mы�s=k�D�R-S&�\�T����'w��k6�Vwm�5�U��[_�b�o��ڕ'[��c`G���t�#TR��}��������ܾy��v�=��7��}j�F��ͦ���9�{<�ǒ����R�9[~ֶ�Y1��6�B�f�蜅��M�ȯ�6;�h������L��[4/0��#��>�}�k�����!��lV!� L������:�u��5���F��L'c S`��ջ��bL�
�.��ڔ89$*���Rc{'\yە��^�e�����N����0?����g���/��h���谉WV SȐjd�kJy�������=*?~����J��z)P�٪ B�Cc"݀�Cꘌ3ֺ=$���Tw��Tq2;Ȗ`,�
�x_V����,�ߘ���d20U%��J�I�	���&��_�y���R2%�����.�x��!@0R�x�֕�����Y�ע|�(%��U
�'�I6W$/�����x�YO<S��K�՗�=cf�$��DF�Q1� :UC�
xz$���G��g*�}�^팧=�A0a(]|�r��	���0��!�2M�?�S���{�	�d�8d(&�I���tp���K�yi��P!Q����4��6�gY���68�S	`�;��)��`�*��9e�������`��.��+ۛ��	P&Lp���� ������¼�]yE���c�j�؍7�����j$f��!�7���z�m[�+�^ xJ߼�4�i�<l�=ýj��VVVT�0Ӆ� ��*8�,#W��ؓ�}�,�^��)�	�*�S�2�lN@"���k�����fa)�$��3�b��X�.��os�TN,�7�Iu�{[0�Z�ś{�����U����WBeK��K����\U�{���Ah\\
�F(��� z V0[u�����	�����o��~��j�}�5��鬒�,dg�0M���n���������ݟ�xS#���������%��3µE !��X�ɾ�~Ϲ!U*էh�(z�,W\���o�\��Ȕ���5�~�y.$/��E�IN}څ;�<�"�Z�KD���u�����B�R�4���z� x�xG�HQ逤-U=E�b��V��0c{�./�Z��*�į�F��5! z��P@���L�Ϫ��g�χ��&�)'����48���@Y��� �q]I�Q��2��X��!�~���1�A�������W�� �Ǔ,��Tp���X���A�ɰ����a���tª*�*��=ܿh69��Fe/�����o�w��J;��� t�|H
;��H�;�̞�`v�m_��������_a�檍1-�ղV�e���� ����;������ ju��(ȔK`����X��g"�������    IDAT��ld�Fe�j�.߬�Ͻ����{�mt4"E9�WII�'����L���Eb�CHFm6��}����_��z��yj���m\��-,�#�g��"���:�iŊ���m묯z�2���i݁���K�W�sj��+�S��V��׭��E3 2@Ϳ�hU�"���;M��,�=�����j\y.�]9��}�^��Gv��GW`�S|6���[����j���Y焫�1�!?���l�q1/�&0��R��������_~��O;6�#�j�"�mF��cV�D3j���FR���������R�����`��ӫ�$*1�#�bh$c�Y�g��I�9�I���iľ�~U��,�})���;XR�Zq���׌d�H�X��&"\s �^������ˢ�|8������%ߟB��/%�.w����&��=ތ`9 ��H���j���G��N��?K�W�SD���=�����G'`��Ɠ�bBV^\?��wH��^i=)qIgA12U�s�r�n�L�PH�l��c�b_�$:1,Q���?���_ܱ0�?��!�CK�xj���3X«�S�P�[t0�K�t�1h�b�F%��H�tx4�k��X��Ѣ����
��2/T�:�\����������ؖ ���}P%���-�!���h��II��S���-���ޏ�7�ʍ�0��qm�3Y�Xcf��4^U�ԙ]�ʀ��|x�g��^�̭1�Y}8��8�tn�&@�~9H:���j9��:�Ǔ�}WJ�J�|�3!	�WI�1R.�^�cbS�r�� :9�����PP8�N��I1��]�&���Iy�/'}ԯ��W=��ɺ��d����P�n8��-��9ю�F<�
��1�6T�s�C
��5�X	���&��X�vh�~�����ͮ�2[Co���Xo���q��]����}v�g��ط��ؼ޳	d\4�iY��aO׽K�!FOb�.�{5�'�$-�5+�/�g~����v&�O���r�"�TRW� ܄�)'�"
2 �J�.)����y%����u��j=)PY��z됃�L��n&��#�"��=�����s��
jl���)+H~���J��� ��4[�g�k�����b��K�u�8��G�|�i�EĂf���ݵeܭt�n���؁�Ϯ�
ô ��k��M����ơ�A��3��)��X��P��ˣ[�Q���kvU��G!/����H��X�"aHɘ�W��Q1� �z4��-�Ci�3�FC���1��b�o���~���G������]a])# 8d���U_������������}��A�q [V�Z�h���8��$���ҧW[P���ɷy��s=���Ӟzx= 3C`�Hs5g��5�O��Z�6�3�5��_x���-7ى6>��x���?�g�bWJ�����]u�y�O���>y����y{�쑝ߟ�`�+�9L�@:{���Ѷ��r5"�i�l�Ԗ��WYi��"J=a]t�uJyi~tG��Fc��A�����)M�u�����`:0����1��9�]���b:��؁����c����B�;�/�e���s�Ě
�GA6+>֬�� ד+�d����lQ��4?��O}�~���lR^�l4�L��!�
�	*�3�P�����'^�ȍ'�o�L"͠�a��᠚*�~�L�"��W�`�Js�$qm��<�2h^2�9K����-*i�;8O��������C���y��%#e�Ag	�;�Ĥx��!_w7]r�Sr�k�!L���1I_����� ����^;D`�� ?�^�3�W��|x,%��ٳ��r]`-U�ڱ /t��&������;�@CI�g�KՁev�=���n,u>��(�aǞBO��Kk�%�!O�Z����:�&Z2���S���S�F;"�a�NP=Db��JH����|d�����=�E���u SVP�G���ñ��lt8 x\;y�VϜ�E�N�@T9(M�vX�'3��[�No�6��uOn�u[r�E�����"Kp�P1�.�c: 0mc�u�Ii%~��R���G4��c;*'�z>3�D��4�H�˝���Ӯ5{�Ui5�6|*v0b�'8d��� �Z5]�5�g�����Ȥ��'����@���Nf$V���l�Ύ�QU�MP�ZpJT�0�k,z�$%_�#�s�Ӎ8��%P��@DS,
��'�na��6&�jFt�@[ģ��b�5�þP%��� ���}tH�$�A���=΅ę5�_���	n�爳��06M6��l2��o�i�Nt'����w��&{�M�����ii� ����h��{fw�����־q���3�Y�{�Gs�7�VGl`u�Q�FN�A0�U5u�	�*șe��T�.�\a���=��X?�����=�:����tj��bLCف�)�#T��O+.��s�)��-G�������ܷ��$�뚍>������g2[0���4������F PF�J(V����˰y�yX��-F3.Ɓwԡ	Z%%^��"�BL��wHYAlԭ���*+?�@b���d^w -3C��>�$����CE.�~v=��|,�z�"���Ahs}D����m6��P��&21T~|�l^��x)wZr�����������܍���QULε�D��s kc>��dl�a�f�[L���+��x����W�u�7�[��=J� ;������S��?��>y�]v�e�=e�Z���hru_=ߔ�䢐���修�G�4%�S�z�<2z���WLĞ��F�b�&֪��3?��X���?g?���l����Rz���A���w�-�Ky}&S�(90E��{�sdv�W�O��{�C�p8�Ѭeռm�x�h���B���;+��R��}��
�1��d��e\;}0�u��`zз���(�Ǵsj۬��d 􈎧Sy �ha����T�t�S�b��f���!c#�>q>�20�tm��GS�N�7� �0|DŔ
0�o܇L<1;�́���iO9��?�b�@��������U����k���jVou�ß�'3Y�3a���(0gr �Le|�J��q`��H�ʕ�^�b����ɈHң�����Š����6�ܟ̲j�E�nC �M��,�!�E?�';�xp~͊�^_�dc^UH[��e&'N��m��1,��������VU�dRI���Y�avm��;�(�����A�O�Ga�8�}�8\�-IY��]�N���zg��v��5+�r���f=)�$�pp�����*�y������uuO (�
 ?� ��ȿ�	,�zGs0T��:|Vƚ��`�S�����
f�n�5K-֩z)��hi�b�\� �ӊV�\7��d��k5��3^��vp��Â	S؆7P��6m���f��ɳ�=�HhP�p`:<$)��-��(~�͏�L��Vۨ"0�o��Vg��t�0�F����� f�5��#�=��3�v��HL�J)/��H�����a.�C�l9�q��:�b��P�E`
�L%{2�bɩ7H;�*�ޔ7��ҝ��z����i��}>��ǉ��U :UC����8�K������"�#��9��ƽ����|ܰ�8d*�0�Ӆd���_	E�����zEWCT�U�R_r|.U��*��3g��H��cM���ّ?�w$���zg��#�D�E�W���6X����y��հo��E��T�����=?�*{�55l-���]&9���ѳs��3wح���=�[٨�j�^�Z{�& 7x���d��A�|]��]5��s�i=�^�5X��z~�DP}�˿�=��E���^>Jp��N���+��p	����n�b�;b��+��dʡD�Y�����j��M���`�J�d�J �q�pB��j(�'ך���0At�PSV�>�V����s���R���)��zh:��bꥹX�$p�k�j�bB�T�<�2�ku ��r�VǸ	��F�]����~�نx�3�s=çïQm�1�Zϑ��	�8UI�O�'�&)i��H��39���y�jw��[yEUJ@�l���li�z~��+����s�;�o�9|��V���T5q'_n$E1Zel�����=�v����~��7ڇ�-v�K���A��y��� ,���}����}�����GV�7l��q7; ���6}ܙT])u"y[����Q˃�t2|R�{��N+ȇ����td������^����������k�)]V�C�ufF�$ŝ2�G4�M��K`Z���rO�x�,�U��Tf���3�������Y{vwdêaSk��Z����<ϑ=��<rx#.8.@.zLQmM+W��]�D`��=XE�̏X1\Le~���A�0ق�����؆�+�d�O��<t>5(��z��r八�xL2�H�vۚ��"��,S_�1�9�Dt�!s�	����Xs:��袽�%g�7�#vݶ�3b�6�/�"�5������}�3�`�;�r8 ��k�)�0�C0P���������$�ɟ[
G"��#t����`�+<��h#{r��`!�d��:N���rjH*�ur���_5�UP�h� � ���{�
	�_���}����㈵R�� �EE�1�8��sE)�6��[�+`�tʅ6z#Y��Ty �;���=��"�b��,�J:E`%�� &��:���f?$q�x�t��S�T�{��l]��] �!�UP�D����L���G$+1!���\��da�$����i#�3�5*���-I_\�BS�T�R�JgM�m���1����3��'D�!��و�^�FƋ@{�`�T���`�
%�4�N(�R���5$����+���`U�Z�71�r&�/#����U��z�j]k� SU��S�D��`̆�Q�����	['0��=�6bd������4�Z��*� �0ju���F`�9��UlE<�H0��3��C�{����֛�!E
V�	Rވy�0g����Zɿb�5��q�R^��a��ݶi�Qɑ�jpݞ��«�An1J�É͆��y5�H��R����B�r�f�vM�9�	ǀDT�� gU�]9#Q��S���E8��� !Ef�I���,;v��g�.��|	i�ZNt-��{Nq�d���"��Q-S��Nf��!z�)�U�D/���cw�
���\�� �z<�.��l���m�T��������ֶO�AR��_:A���f��7��?�k����sS[����X�	���:��Jq�����\'�\/�g�P��,cm`�g�^�^%j$I��V�-�e?����8�\��>Ql(H���R�	>_�x�q�I���@5���H�a��\C��l�ʦÁUC%��ш�9Z-̀���bV��<�<�U�Y�Ӵ���]y�)��X�N�aݎ~�ݨ[�۶N�jUZp���
�*-���J|U���X�)⇲u�U�L&�G�Fy���/T�=����]{�܎���pPY���(.vͶ;���l1�M�uwm6�,���4�D����H�&χ���̿�/DUoe�r[�����h��g>ᯭx�H^?��(���R��	b,����8�$��Xv�����ne�)>�7�	��=B��d6��U�#���C{�u�����c?y�sl���Sv��51�q�nd��/���o���}�o�چY� �|��8w��LWbWo��ׯ�;��D;� �Z-#ex��iu2�	��ZO�ec[oWֳ��|���?�3��kW�ow:�=\C`|-{,G��?����\�ł��"��q&`�����ؚ�}���c�������l�`j�
&A��D^ذ)�������n���fU�a\�g�#O�a��Lt��u`�3@mq8��h@�?�� ��V�w�=5h����4a�d��m�ݲ�?��ᡍ�6W4j
�Z9[[r\�J*:�Gu�g�1�lgצ�	�M(gt�U��D�ѫ�9����6,�� ���LhTkOv��.��O>d���;̏fULw���_���۫��UU�¡�� ��d�|ni�}��h˗*�`�9��ј���K�fs�G�T�q ����^��������4ʁQ�a D�A@$X9��KrPiR�F		��`x6�䓔��y/B���~�#R2� �U@,�YӇ�KDPE�2�ju:��#S�G&>zT1GO���Q��J$@^FIl=9!h4�"U�\�eLEITK�p��u�f*[(�Y�˟8�հ&.�,4𽸷�R��^�4F�\Z)?E� ��J�QrrE�U��6�͹4Q�C���~�zfļf�f�py�_�� ���S���gz�0g�I�O7�r 	�,�%�M���*�C|~]ɟ9�{0u��2	�r�K@N�a��!v>���6�����S���.Wí��2����U��F�j^10��� dh~,�S��u� o ��YU SH��Ks`��}��[�m��u�ڤ�Ί��)4'3�V�6��68w�� � �>�2��J<j��v/���:V�R�&��ª���[6��f�uY5E/.g����T+���p��[[�6� Hz�sf�ӷ��`�~AW[� �k۝h��U|�]ʶ��~�2�N3�c��}���[$�I�^��H�[�/��DTU�\��~��k����o6��������A�I�T��q��#7oH`�ϖt���]1�P���}���P�xI�ڴ��dG���_�b��÷�{o��N�8��Ϣ
��Hv̆3����g����쯿��M�k6o��B��ڼ���H����w�O|.����1QA`U	��Q{�z
ɬ���s�9w��-�K�k�I��<c��D����5�.�^ <F�=��"oq?*T8�c�>+�hj8�Q} ��'kbc*�����Y�ӱ-�#�W#��x&k�]�:�F𹽹n'7�l�Ć��>i��ٶ���v�Ԧ]q����4�մ�\XVTScM��*U����?H^��=2Q?�-�������߰���<�=����q�}��cO����#�����F������O6F��f�\V_����(����R.�v��Ls�w��b�*�R����X�j����r��"�E�ϖ�0o;p�y#	=�'f�'gp=��u�ee)�h�~ոXѤ�Z�T�W1��O��=��w�>ٷ학���n?����+� ��*d���a��}������K����i�5z'm�)T��t�
�c�z����9S�g��C�K��{�`�Հ����U�qHm�&H�5�oZ[s�o7�p��g?���W�J+϶�t9�]
ї�i�c�TQ�zn����W���Y�����=�?����=�=g����BIж]xU��ϼU!L�|c�PO�`n<_XըY�$zL���3�&�E*B`2
s��ȕ&��G6!0�T�@�$S�P�+�s����̆�LG���[m���"'�,zUxϐ�`*ڜFG};��\�G��6W�fP�%`�Y��x��8��3�: jUq\L�ڳ�_r��ٯ}؞����ȁ����l����lұL8�]�e����H��Ť�s�����Td��y�J0�tb�ȍ�J��C[$��g@e~I_�Mx�����@j�)�VU�d��0O��R#+9m\�y��-�!��P`Փ�ҿ+Ⱦy����	�Ԩ�1aU���2������ԊM����j�	z�A���$Q���b�i��6e�bv˵��*./��0U5��!/�=�`Ð𾺬��n
浲�J�萯uWWx! 
���@ep��DV[���a2R�s�����ȍ�DTd	y��Q�"3��*����~���u[��;���&�.��y�'V \�G�^��� �@��cܽ6L r��|k=p�Ic�����޲:�x^�"�N����%;?�X7g��S�b��ya���~^�v�,b�P����뉥w�q~'��z�K�L��ABL�N���&���1%"ã�zL�N���TquG^J��(��Қ����0����`:0m0%���*�3=8��y��"!����m�Xq_xb���yT��(V��ٕ$���ʁE�l    IDAT�	R�c�væM#kʪ|ar�"lX}�%�'�S[��C�y��+� �Z�K�P�`�At�kI�P�d��D_�����G��T�G���ę�_T����:��^����� ��1N�T	�����Z���\8}'R�p��<b��_R�XLM�-��@]��!e���=��{I�J�9::���o�ɾ���+y��ī��M�>�j�H����;������K�����b��5���"��"1Wb�*&��}���#��*�%(���R�:\�c��cy�莫�/��Y
1_�"W���C���`h�*�*\��s�㣈F)"��S���J)I��>� t�m:��� ������a��敵kS�\��e�7��.������������m���,Ӑ�u�K"e�k$��-�IJ�w�<O�%.��+=�p������*n��e��8^��Q� �k�-l8�A��p4��þ��ڳgw�������y�=�̮��3k�Wl0F_�jͶ��p�����B�x��k��0�M����$�Ǜ0�R#Е+���P�-	(�}��h��c
��V�{�y=Gϖ�SZ��X�KA��R~N5����!���_�J���0.j:ر����5/�_|�[�/9m+�z���ta�����g����_������°e��+�Zx_1�W�	���@V��$�\6�<>���燮!H�H��k,D��۬�N��Y�6���Ȯ�b��s��o���:��r�A��*����-?���|:q�w"��V��	Ⱦ���p����;5�p�s�s	�7@�4��ս�:I�_w��;��mR����I�8��J�Hh���p�m!W:ش?��hb�)*�UL���� C"~aU�ق?����
�zÑ��k��3�S �͏���#�jfk+����V0_�CƌZ@˚+b�8i�Z�T���$��B��a�t�����d�R��k��~`z��~��`���a�/V��U���6X*�����H���v��*!̇�@0'D�:LB��OÒ<ST�O�A��:! !�&��:8�,D@� p���|6��e��آa�x`-������T�;�(��7{%6�`��H�yb�F�8[��	�����^�ٔs���Ԑ?h����]��'9�I:�,�5f`��eJ��a��b�Q�?�?U��D
+%�`l�׳#�O�3s`���)���ZX��&t����m(�b�	~7m}s+5�Kr�J�l1��c����!����W�����y�CT$�0c�KLHh�3͉MT�=��y��{e�����0�P� @��b�T����<��UQ1���e��~�W���t��`�ul�_(邭��rg��&=]k�W��\� ��T��t����\�d���*ߋ ��Q�^�'^&֒�boF�B���f��+	��r/����M����G68�3(��ܴ��'���CȘ���mᎍ+������k-�8�*� Ƭ����*�rT	L���Xk:�n�IEDT�B]EB��9���ȧT1#��j&4>��{�D��S����Y��n��]� XIt���� 5�W�c���uj� ��	P+�n���$D��+i�}s�PF�U�:ֻ��K��JCΜ���gL=9**�u�9�tY�o/��pc�"���V|o6�I1 �d>��c@���>�ۂ-��	�䨚�:���0gqfޓ� �PU0�kѳ��k'�;����@��M��6ڿ`�ɾ��K��_���M/��*�*�iT��T���`�ñٟ�v���'�l���l�XQ��ֶv�#GIoF%����HÑ;U�ٯU	�<�5!�� �^�I�,��ZП�
&�9��[)^gI��A9���㔳�$��]�&�S�o  C��9��59�".�,�(����C5�|<��p���t4�Y5�V���=����N��W��+O����=���-;��a�O�����(��Q}&���f(ֵ�~����0h3r��2F�_�t7�մ�QR;��)���!B�⸌u{!):�c`����C�����vq�O��>n�>��=un�vaj�s�ն��6�5� �գ��E�m�E R�[-N�� '���f��}�T�9(�5���.U����EI�I���6L���С=G���aį�ʧY����Nb�qz�l��	>�����c�Vv�w��}�ؑ����/}�g�m7_��SO�X2	/�����[o���?�+�Ї�v��5�0F�e��� PQ
P;���I�U߽��Uv�3��>��AiJམO��Zؼ:��|`[݅��?j���7؋�[���2D��bȱ����Fmp�4�0��ݦ�J�������Oۭ�}���q�:6�@9ץ�=�gȭQ�T�*�h)�
��2�w�+��67�{b�*<�$b�<��B`
"`{�?�j8����L��ۜB@`��i	h��{�F�M���4�j\q�zCsŴ�Y�&&���ڥ��`:ˤ	���i�7#UL����1W�#I����TTL�#ӛo��~���=o����V��bR7�87����v����y�3x`%��/�w"x�d1WLi �ڶ( .r�v��]sf+�Au5ث���g�b�y�?CNT���%%�4��]��\��:�ǹM�C����Sk��뮰+/�ܞ>`O>}��~��m�u��o{����W�|��������n��v�P�M���<��8a��Ii�(x:��N%+�,�#������5kb�����]�Fw���7+��ʪ��&*����x�mZ�X��f���ם��qV���78�g��L�R�{I���N�ɐN�p�\L�6���!�b��C��Uk�6���H� ��ͦ#���6y?��b�^�ٱn���j�ˍ�O���,�zJ��D�P�T[dTOER XA�0���H	P�l �Ƚ�r$���2`Ӱ��/�O���H��i��0�{�**znK�}��2Qm2��ԩ@��mp�oG�����y����VNX�����oaM�(��mx�ǾCV��M�lX��J��2&$d� J�* ��m�d�g,J\�QPiVjTѕmANLب��B�&W\7	 u�uV�&�!����b�qf[��6�ϧY��P#	�SB���������TŴ�'�[���	�Ƣfmp���6��k�!��(d>
" �[ޟWT!}4I7J�\"D�W�̈o|���|��
�#$^��-`�p�5��%+� ��;�B���^옚�@b��?"@EЏ��"�`�s�D���K:���p=R?,�WC��+d�Y^V9c����9	ON��R�)�w~��]�`fs8~g�Es&�h��r�SUD�S��"�$7��:í�2'&3�u&(�d	��m!�ad���̪�M��Y{�c?����?��-���W���N`��%���pj��SSJ̾t��v�`f�ƆMm��:j3a��d��SC�M��	�F	F��ɴ/!EJ��f��l˼~|�%����9B��1�2�s�S��y�R%�ɮ^8�*��v��ccֲ�y�w�\Uc�LF�3�<��U�C�e� y�����=�l{öO��5W�����:{�M/���-�OT�K���{$��˰�#�K���5��3	�D�yXT���$r&L��}� ��@k'� km�g+�,ɠ� E���;��*>�`d�����|�){�'큇������6#6#?X��:d�"M�m�Y]k����:�B��^=&��B_/���9!)%a᪬$�����?���y��e*�S��1"~��K�4�Z?AJeB��J�Ql^p��UO�s���Շ�l��C+��=o�Ѿ�ǻv剎���o�������5VOI���8��;8=�̾��g����mv��m\���gP�	�C�F�\�|$r3"�r�(����e��BJ����˃�%��-�Qs�W�6�6��U[{Ǜ^my�[m{�&�X����'�g��2�[�n�z��㸝��Ρ���}�>�ٯ�J����*�irW�
�CH��x�w����LjU|����S䞵��N��TL'(8���2E�MDp��.Cn���~���\y�b�Lh�&�����lj�hI@u}� �k�m������E� z��V�m�b�G���H>6� Na|P���R1F��)����G���X��ڳ��2�g��!{�ɿC�;���S����n���|��4^1�a����O�H8!}����<�]�My���I`1�)IƢ���#z�-ņ�����w�7Ts� O@�J艕O�3S��}k��^�k�#�{��ȋ7y��̾x���ͯ����o��_�Fƚ���u���ڿ��O��Oټ�f� [��v!�(��oȉqat��U�}[o���Wm�+ox�]���m}u�C�iL�hڃO\�O��E���g���엾����gϽ��]y�6?�ɇ�8k��[v����ĺ��[�I�*�HR���g}8%�Q_t9���������fmuj�b�g7\���3���a�����`l���}�އ�;=m�z��6���Fۮ8�iW_~�Nl�����Sg��g�sfn�w�j �9{0�!��h�F�L)�B��]�I��B2=��`
��Y�]��0�h[�ճf�� 9��k���.j J��g��}B2 ��P@t���j*i+�8$+��$[!���qߎ����t`�^y�N�\�+/���F0����=��E��?�vgÎ�^��{��\oٙ�M봚�з�{��?��hj�EӚ�MktzVo�^�M�⃙����%&�.Ǔ�@)@d ��:*7��T��@i��Y��`D`:�k�)�Ŭ�ޒAPM=��T(�DUJyǕ�� �����`z�z��6(%f��=�;�f��*��{֚.�b��Pܹ*j"#�0��9���kQ����_����G��U!�K��:-�� � �4}���D�U2wŔ�J�QJw)�A��� ���F2Ğ�|h�Z��}5���]v1���-�$.�
�D2�$�5�wS�ҥ�H2�CT_��C2�$8B��!������ֽO�*��Kix$mو����q��AtF�PV�܋��^!��c�]��s�	A,��UP��g�WGV��S��}�^g|�k��Ӓ�X��+��aVx�l�o��=n��W��>cG��u6=�i"�ʾ>�)p�fVA8�"��%��e_`�^��rn9������ɨ�~�V� ."�q����L�1�x��5V��&���F+������y�J�-����Y$�P� ��C�m4ط�ld�M��lۉՖ]vrͮ�┽��W��{�=���mm��W���O�L���Q$۽�D�������׺�_�o|	�1�%��A���u�뗈��{�DЬ�-����6���B>�)Q	E���E6�_l��n�+����s45{♅}����7�~����#��7�����.I(�*p0o���q��5AX��^��"����ȋ`Ҍ.���,"Z��"�%�,��z����X{�����J:�/�lΉ�y�+B�*�4���ƺD]���+���P�Bwa^ٰ�Oc��p�V�#{��>�޷�^}-G� kR�T��1�x�0��q�}�>�o��D���ح���g�jQR�-k2պ/��z��'u�;	8	+��et�C�ܷ6d�ա�f���믴[�x������5�����޲�Hz*^�W�d����aeva��'�ݱ�{����{�G��s�c/0���+T�hc�f���znq>�IT��p�%bU�k�Xf����<i��U������<�~5^�l�g��v��:����h�Þ��s
�O�7b\�l0{�����T�MC�r\���-��\����U%p���l�Ӷ6r�����G6���{x��*k|��ߚ�	)$�4z	CA@TPQqt��q�3�et��mD@P�"�[�I� )��'���������s�	�?_�]�������<��k�֎!��<��T���np9��\�R��9�J����=����qX�_p�m�[�
B8P��cx��>�ZIy �FE:d��8Z�*�Ƈ0iΐQ>,ѻ���wp��V��V��-��j��d�:�+j@T��(�����	�P����4bɜt�X-V�*�QL��[��I,_���M���S�"Ԭ�����dR�,��
���/n{�:g%ŉND�FCu�Oi$�S�c	E�QAy| ��N;n>r	���R��+?��~y�x���1�-�����8�I2pY��Ϫa��¯�|Ϭ{�H�x�tV˧6�H*�Rm�A��������W����/�=��;�x���W-�%����M@Z���� �ۀBxq�~������b�t�����p̒�q��,�qe�:�}�^xu3�|~#�lB#�E<�!T��7+z�V���cB��k���"3"k�R�Yҷ��.&�J�B�י�%P,�Mt K"�!㑈 �f�4��uHʵDъ�Pf �׊f&"+��#����=V:�0��k�V�7y��hW�n�1�8�%8���>�Y�"����_��^�R�V>-̟Յk��"6-�ޮ����ױo���}#x~��x~����6�TG�̭b�T�g:�\n���>I�t��[윫�c_%�<F�+�h6%�>�f�(�-Ho\>H)��0m"���S:��x����8�JǴ�*����L��ۡHV]e(0e졦X�)5����E��&�͙T�d�"�ar53��(��:�F�T������8zT��)�ZK�7�w�o�2�2)�Oj`�\�mxtk.3VU�U�R{��Q��H��.�}M�<(�3�̕��*]��<eN5�����HA`*����ӭK5?���!p��\��Zc�9
�\Q���8{:�w'Js$�#u]n}2
�MX���k:��=�&��6S�2�8���0Բ V/��]E�����i\~��x�Yѝ�d�d]���+�# ƀ�~>�
��Q�Q#C��2��$�Cd�����C*�����1��x�/{>��������j|��+8��H��:�����\�����n�>�KqǨ���4ѐ�3�#R�bA&*I�J�*�AԫbbԨ��lQ��!o`ƴN,_2ǭ\�y��b֔^L�I�3gzP�|u��+�(���q�٨����Z���x#��˕Nc�N=�J}�/P�VQ��|�Bg]�����k�<wH��~v��~.���G"�./6A�|���ѝGkA�]XX��Z(�E!k��4X	L��T����ާ������_��l���1<ZC��o�t_�x���v�O2!NJ���&�:��4�@I�%c�4���&�.5����h����i�+2�b.��y�fq�́S�����7�u����gg��ɖ��d �s�U���N����ѨoE���+/��'-BOF�S�S�,֊��;���������p�P��[���H\��ԕ/�%���Tqr ���v-c�����l2���+-��2�FА�YA�UA�YB:Z�aS:q��^�\2��¼ç"�K�[���p{���hغ�[����7���m�00����M�u9V'D}~��8U ^N7ig�c���%������5ՙ�,@gzzI�D��܉�Z�H�Ŕbu�mdB�c�B�PA�P����P:�XO��/�������y�FL6E6�|�M�Z��&���Y�̰[J���!�j�ĳ�k el���I����wvL�O��n���u�$�`̵�k����	M�kU�%Ī�8m�\���pX�_L���O��l��qw���<��6�F���v����3s�M��N�RI�c1/�"b\�6�@j6{�����B�o��撰8ڠ�AR�ԸƤ.V�	�Lͫ��/V�ֶ�زm?*u��:�t6�Ъ�b�T��[��Ԝ���m��Wvぇ�����3�"K���A��+xcw����0R�@��D,�@���.X+�KuX挪�6�c+�^E�|�����_v�=j�X�lG�9��G7E�޽�m���Q�r���1V9.v%(�ۨ�C�¶~�n��n���.�S�
�xhѸ��Յ��w�p    IDATH�A����K��Mէr�$���d��A�U|�+�s�+��+j�6�5y��1�����ƶ;��/\�U�M�I1� �mQ�D;����Q���?��w"��F8�5ڴ%~���͹RL�:LZ՜֧p
]�Q��ۜ��8��eX�h.bQ�r��j-���}� ~��W�@Z: %@ڿ��0��ET�C�=�ǭ8
��MEQ���^��e'J-
F����"�P>��)�Z�j�ј�4ڵ"
�;�x�$\u�{p�1s0!g�>��܆�}���<���o��eKq��q�e�H���Rx� =����F��;zѢ��Ss���"3��?3���d�%+0iMH)(e҇c��r�f�28���3��ر`ʎ鈣�Uc:��R䩫V-���	5֨�QC�Q`�D�f����4#j�� ��똅�t�1��P�9a���$ƒ_��+�xe^�b1��M=��" 31����R���i�Ҡy�7�\��h�B��X�-\{f��=��jȎC^���9�"u����h�|AM�<��s$�H��k}ʭ}����ّ��\�L���bUmc�B�3O�o@s���q��#��59ڽѓ#إ��f��C)|;,���v(����@V��sč^9���s��]]�ej�xʌl�=��f��H�Gp������S����od;Yᖇ�u�j-`s_w�����&�W�]��8B,�EH�U� ���&<��f�gtu�������}��i���j��ZT���X�ϵ�i�t�����mX�4�L؃q?^i���k2/�h)EiB���΢6�T�+e�8!�G��G�QB�VD$�Dg.��K��ԓ��ؕ1w�DL��7�l��)���{:4����4ݦ�$�7ו���)�N�ηZ$��R���(��܅�[�c���kɗ�R�g�����t�I�	
A�R�y�XL��p�֎�qDBa"�L:��}�$r��:2�X:l�̜>ӧMB&��a-F�������_�~"�
NN�g�|��pM˺փ�3Wڵ��W7��SϮ�K����P�
ǧE�Q�G4Au�D
�\'��"	2�lԅ�$�ж�\�8f��\�m�������?��5U3H��ˇF� #�"�_��h�B���+����r�\���I�4tDo�3L���K45R&#�ڭb?����9W^�L����f����<�,�����Ol�-�}���#���p<��cjB�sȵ���[�-4��}��
- �����a����u�m���yEK	F2�v�&�_X|F&�����9G̞�c����.�%g4FId������[[�cǮ��sC�T�+�}���x���������+�	NP�]�P&��7���U@�B�ɕ��<�,3�dI��%yY\!d�!D�c�����g�DO�t�37NG��z53d��EБH ��4j���Iyg���n)g�
�p�H��s�U�����`�]yShZўkEJfZ++��(R�a�&L�ZȄb�a�Z:]��,N
��0Ďi!������̫�P��Y���W�ąg��ӣHZ�M�Ky�Gq��N��jg�!�x�5�k(�)=ɮ�U׃���n�|b;�{-v�B�VA��G,\��?z!��է"-ء��
��߉��٫/��&��
@oWJn�0���c�j���"I}��j�θ��5P:*�DԪ(���\��7�{O���8���H��V9R��op�������:���� Ϙ�9|�&���#��wc۾��^Y��9־�~��\��#����B-#s��5�ƆPه�x_��O��Gʮ��C꽮hs$i��������_trdX�����K�4"a����۱y�(Z�"O2ܥ�����f�ز�C@R��Z,�Ӄ�>v1�>"%�iw��ă7�� � ��9<��f�7Q��S��8�̟�O|�\��r�h{����k���ǰs��r��M6O��̺�V,nâ#�b�Y/�����F�TF�j�+��e�,G'y5Mg��~�#��Ɓ�G0cZ��w��Df)���:GE�����p���p)�F�t��\���* ��V���\b#B���U��V�9� ��	�n��k���TA)���r��Q�r/R�9q�9��
0e��ɽ�6Ek+J`�ęW̢�I��@�7�V��	�����Ό8�E�c�EPɣ24f�b��K0��!Yö�d,���>���5��r{�3c�y�Y�̤��*��Ag���A(g�E8N��ak�Fe�U��ΦFP�y�n��S�Ы�[���w�cj SX. �:��}��7��h��x���)��+��p6�\����x*�T�>�8�w�:�@���n��Y�=`awI�W�?�;��q�Z��:*Íw�y� �m�$S�ܐeO��]5�U$O454��� �ǚ��:gG�l�YqO�0�urp�����[��7���B8�!�<�vOx��	��2;�����c�[=|���+����u��g�C�J��qk�Oh�b��B��5� �q`�����#`���3m���#�B-��M��QA�0�z~�J�v�X��Iy�l�t�r�\�󏘂�n�+�9��&��ߟ:���%�b���Y��*P(����mxg�.�ع��"J�*b��:g�hT@�`Z4�J�c�:/�HT�����u�慫��W�s���T�bRA0�p�م��	d�xLƷ�tuu`�䉘6yfΘ��&ʸ���z���f��I�U��L������:7����������r��,&�9_��c��[�싯b���88T�h�c5ح�ټ�L�&"�N+�#�K�d��c�֎�>ez��\N�}���3z���	�c��t�[1�s��*��ܬC+Q�3�
���dֱYZ~W�"�̖4�m`W�k��_A���<C����'/ǲ#'##cW�˪����Za�f������݁�LO�'Q2ƴc�F�y5L;���������s]J|������'��­��e$I>���d>F�Ҫ�1�n �:��Sdf�{�C��V�B�NyP�P��`1�v4���jg_���G��[g�KQ�{�y��h����e6��q�`�)���"�;#�cJ�'�IS�cZ�B�tLy�3�uw��&�����:�#�B%0-��V���j�1eh�"%tD���SeA+N��?ՊtL�1�5�PD*/-���S�C:�)5P*ESF)Jո�h�W7*ou�/���p)fu���i�4�}����;P��Л���W�Ⳗ`),�e�+6[�qW�y�1��X�����-x�?��4�?]@�iN�
�Ԧ��0~��?��-�䡕��H'��ϯ}�6q(���o��t�~�b>�;���W����FB��g>�	5��9|���������T�"�&��t4�S�H6��Q݋��t↯��N�*_{����a�֙�`⤌$5����w���s�f�6:Z���8�GG���YSdV� ,^���=��_܆hj�қ���	�H�;��Ѱ惀i�hB��ʜRW�4�A~p&����?~
篞/����q����ݡ�����ad,��s{�4���CC�ǣ��%�I��m�ڎb���W���^C��*���jKM��TIu4���)�e�^������5����BOHp���_7��ZC�6���|��wc��Q�����+_�$V�E�\2Y x��!��Wb�@�M�"�'S:\\v��I���Q��b1ޢ�q!V���8�����k? ��0�mͨ_|F�\��^�Fi+3�n|�S�< H���"xm��~��{*��1�%X\��Pm�_�ר�8�{���jҠ���$A[�)�h�T�LJ�f�|�;����%ň���i^"B���I=�d�nU�)-�U�-nuF�eǴ��Zu�j�?�to�hL�0J���QeAg3
�Q1?��kǔN����P�$xJ�q�1�Q�d��H�c��K�]��/�V��T4�nƭ�P�H4��3WQ��kj�Osk����/�פ[/d�YK���Y�A��L\U-���u����<Z���Pk,�����߽�%cj��q���ˏf��o�=����G9GH�;����hxn��G�����a�q'�v=5���ݡ]� �rM�S����%��-�^ݔ��V���dZx�Y���"��*�A����ۍƁq����翺�G�����A���S�,����k��B�.ͺ�2>MU��W(h� 0�X�9kw���i93�0iEOj�t~���Ǎ摢b ܻ�\�3�D���:�VJ�E�"Ҭ�Y�JO6����`���s��r�S�ˤ��d�x.��ܴ�i��~��N�i�2T�� �`p����Ƌe��+884�]{�c�ރ���/N��+��)G���&&vR�����MT�>J�Q�&���ӎ�� �Z?'{<P\��]Ǝ8�r�ZYL����x'rĥ�YZ��ʹܑN���S1yR/z���ͤ��G�[�+�Ť	ݘ��)�J�X��?�5���[)ߣ7���b�e`�&6l܊��o�[[�aލ|�!�V4�X��L'2�=Hf:�[D�&�/��.���TJi��\⯚)�K*�qL��zvx��N�;6(UUu���G�J�l���!=�7.��F-���~��F.%3�g8��2��"�q��	z��\{��8��%bDp�Ω���O`Ʀ˖��o| Ϯۆ
M85[؀Jaҝ�xq��=Qz�랺�2�eew��a�x�Y�6ׇ㤅G�4����Q0ʆ	���f0��a�\&D��_�tFCa��!_��xƫ��{/���~Z ������M�3)��q�Y� hr����(��c|��6u� ��R�oK�'�h�1VD�^L�� �A���TBdY�!K�ʂ��1��IE� ��m�"�4GS�����#�%c#�)L����T֪U3֋!����2�t��15�'>u)]�P+Ր� �p5�xugs8���/�����n�9L����� ye3��*&w�p��g���0!�ȖU?��[���\[5�p�"�;��>�
�������j��E�mC�'"ln��J�Ώ���KW�XAow���u8��i�5��Ě�4�����3N9�L?�~��_b��I����=&��[�c���~�g7�G-���I�Ɏ6벨�J��}�F��,��+f�_�4�Q��.g�]�7��S�q``ӧNǪ�N��9��m|c+�::1g�4�ۻϿ�2��ưw�N�a|�Kq��ˑ�*�"���/���mE(�+�b����z��mV�͛t	��\�����X&���֗��y��-n����w܅�}�J�����՘ԝ�;Z���b���a�a��n=v�ىG/�����,�4�Ac-��߮�m��E��YI)���~�<]X�B|j4��RG[k���*:b%|����KOBN@��j���Ř!�޾��o��[�}y3j������|\��(�RA����������%�ҽ�-�zPm�vee�q���ŕYa��r~L��'����G���<;Ŋ-��p}�P*��l�<��h��ՆɇY�(�#E`x� �͞��g ��v���������@(كH<"�d��`*�N�jl�T
-\1�~��G �ZX	F��z.���tz��YVԘ�ǐ�K���v�s
�)f�FC%�
���q���ZS\y���Ha�qGN̏ډ�LI�2�t����E�;�zT^�X�>إ�뮎rM5eu흅R�����$hQ��~��ɮ�I��.�7*VP�(�Sȁ�.�q�N�i�����ĢaavNKU���4�`�^�z.�ҡQ�k��+o�%G�!�3ϚC���f\GD^ʪ�Ns�*����G5Z�%��5$��K`��i�_ ��Y�'UmO)�:�8�
��GG+�tO��+�������&�*C��&F5�����*�2�*�@e@�.y�)8���1�K���r&.�6������{��}{����d�R^���4�WA;�L�Uib'p�kk��b��z�C���u +�{�{7�^�f0hd-=W���k u�hmF��V՛�j:@׭v�@2Jx�s9�����*�4Jc��*�;s"�-��%G�����bꤜ�RM�h7���T���A$%�v�i,X���a���(����c߁!���E*D&1G���c���Ğ�R�Ƣ�gFqNּA��Z�R C�)�����K�Δ<��-�`!A�x��1(�5ѡ����I�Js)�6��VJBm�k�L�#�WXJ���fRI�iL�؋�'��S1{�$�WΚ>TW��G��?;G<���CGJ�d��i�oU(����-xᕷ����зw��Y$3݈�;cL ��x�9bf�`H^D&�1�w����<{�^1��{>&E{7s��^��E��:�������z[�+\��+�x,93loJaK;�\}�D��z9�fy��8�N�����EkN��. I�]�;a1�+#���7w��_?���nE#F#�N4H��L>�e�f�����+
���ִ�`8ͩ[��.�t#�����
�ZD�̇o�k�����	�+lɗ�k�����,�ex�_�/���i���T�Ѣ�F]n�8�C�M�b���޴�F��)0m��4��Y�|G�gÊCe\̸���4kk��SiĻ����5*DB�κ�V��24)WQ�ܪ���,�<u��!0�}Z8Q`�P	 �1��)�)����1�͏R	o��Pym�׷���Z�7u���z]�	
LG�c�����"�`���F�%0%�w�͏��Ck_G�^Ǵ�8���\\�z%&�4���kx{�.���+v�<��Ų�NѭUPd*�K����(≸8�ZIߴ��냶*����,F	�j%�D+� ��"�b�Y
+@on���7܍uo�E����(z{��翹
W�2�����
(����_�܇�/8�d52��u ��ތ7�Pe�Ğ�����͏\�!�<:x�ѽ�`Ց���}J:x���b������?�r=�D,��Ka�������B�NG�v������	����q̒�µ��y3��0m ���������9IB�S���|eU@��f0m����$��m��b��vL�����5֜:W:{c�e���G�~V:���z��ﾀi:�<fwq�A����?\�X��T6�Y3'����c�ܩ�HP�ʍ�P��?�/�q��41qbWL�rm�e7'I:j�ՁGT�5�ȅ�����KO`�pTi����� ��S& Mm#�݃U�p�xz����h>�f�2�f)w���X�?����WB;�+������7:���Rɸh{Ĺ��J��ȏ�Y�#ǿ��q�{K��	讑:��q<���(J���58���H��֊���-��ݻ��p ��{Uq�.�I+K����-|������LD,E:��|,aգ�:P�VB�3�&Tz����HTԘ�;��6�38��X��ɘ�l�TA~p�Ѽ̬��t�sj��P��!�u�+���Ryk�C�`�
\$�Tޞ���"�K4Z��au�����:�GipD:��X\�GXhkSi�� J���ӓ@��V\B�"x��sU�@gRu+�r� 	v̸���Τ��¤�*t���K�m���L����JS��4�v(�	�-��gT!9��$?�����tzd5��> �N����s��v�i�m�UR'%#ń9e	4n���+4�릾����wKg��KNR�y��j|m���U��<rg�vL�ٞ�W	w�-�.i���yU�v��(��Q���=)����R�y�L���4J��hv��^mq�{7��Q��� J�j��-2tl�j�6H7FV���4��4�H�HSA	��i�Z��l�y�'�-�%�E�L=�H�pR��)�NYc�h��(J;�>�Q�(�c��-�s�R�h��Gil��ڥtf��5�'��y/�& ��H1�7�Qۥ�    IDAT�H��� WH��+�9Z.�(z�
���{;v� g&W��������s��g�'�р$&�v��q���O-�Y��+�|��2�Nحs�>�9�2ϑ��8�k�L;��0�w{� �:Hǂ{\�K"������<���:bҍ�.����c͙�6Z�g�5�kl�x��X��T���\���{�Z���_�N,�2�g!��3�ӳ��mK�W�B��^:�ց�q�ow/�ی?>��'�[�ӏ6�A,�E���L�DJ�De{
0eǴ�q����~�JdO�ɖ��^q��u��_g��g��C;j:ݾ6h��:��l�ˌq��m=k�̥&F��J-:MTUΎ"Yt��8�-&Gѓj�³���>v>&u8���Y5K���ͻ������Ww	8��g��+�
�����/�'�Ʀ�!�Y���<��h��
�K��z_ě�Z@��
o�|4����֮c)�{! 5`�g3>=��(���/Δͺ���aaI
{
x]��C��pd����(Y�I�d}Q�c�8C����Ɣ�Y"���J�T昖�uI�Rv��t����lt�ǟA`�i6�]w��14�Z�����L�hs,'!�`�q�<����Sy9�� �X��iRr�l��F啑�V��{B��Sv3[Uj�9Ǵ�pq k�����Ř�����v�c����[����j�'����/�E�W�׀i���]�?�����;�P�����'8���]�ۖꄹ�1�w�U'[�'�n�j���v ��LL�2a��KarOu��8v��A�d��*�?�/l�C��@�0�L��+.>_��L����������s���o�C����&�(p1��N��p+v쭢X� �M٨MQtf�n2�vY@�F�U0<���~\z�r|�KE'Ƿ
m��o�����g�/&�=��ӧ����Pȏ�٪ m!�#�h���g��0Ν��E�G����	�v���$����at��l����u#Z5Hh�5�@"
�����m���ǿ|�>_����ҺW��K���^������\�AtfH� �+�}�����)�ʘ;�\r�y�`ͱ�=���,YT��\uݷ�iW��T�3'��'H�Կ�ۏH;`	L9�Uͣ;Q`��KOFƞͦ{���/lܲC*;�^}�w�{�K�0�oࡵoⵍ����Xu�<t2�� 5"��w�0��;���On�x+#b���		�R���F�t�LR i�ڔNy���.�+V��_��[�H~��%|�7��6�^:;;1abb&� 
E�,c�2�8�,�������'c֤t$"�	_��0�n/n��!�	��T���`���ڥ6C��Z�T\�tM�L=hEd'~�D�S�f����Q=͝M����Tj=0��hLC�Ѝ�i�LYֹ��4T��:��2�G���PT����B���Q���<6�<�l!��44���8b͐��*�\h�Ύ��Tg9i|c�eG�}e	�;�吔��LDYHs���}���s�����e��k"&ക��		��U�y�L^-ӱqE֡"Y��C��v�&��v��S�첹DGiz�+��i=\�n���l��$.��{�6��h�^�w�Dg��wSJ�6�'.�p�Ҡ��(!�ˏS-�;0�&Y�wO�Ł��%��%�k56Q{�5(`ۋ���*�M�')�,� T��y���k/��+&"�i�n-�_�
��k������=���2�3C�?̢��П��:�+��ǖj�]�L_�3&�> �*��;�ɍa`WV�n�������Z^���z�@@`�����4d.��@υz�������ZE�UFO.�EGL�E�©���#�$M�h�+{��U�v�u&}u��΄������`�νx{�n��s����Tk�6�3��H	T5��ΤDFlD���8*{�ET3�.��:�ؕFt����K��:ס�A�?�P�K���t��+���rzH��EB�uzl39q��/D�yEM�e4�Um��Q�ՔJ@�
?��!��:�hTT3"��`�ܙX~�<��H̚փ);1�3-Ϗ`�YM9F��#+`1i��'������{u�>����xj�k�܈�;��B<���N���x�8,���k��E+�Ȏw��硚bE��!���N�a�d�0�"�J������8���A��џ]��I6<gkw��x,s��~O&6g�WШ�%e�E�9u1�擗c���ĸ�&.Vj�FS������]x�mh&h�H�׿FE�����Ja����%/� �ZV,�y�毚}?o���;�{����Y�rsI����,sW�5�I���k��K�\g�jn��.�g\���J5��O`��!��Ey���e-KeȬ�Ĝ�%�/�F�N�sYϕ�1O��m��H;�1m��`��/��/S��C�*��{{$G`^L�Z�����l(5ёI GFg����
Li�Dj+G���(�H�����!*}��2/����ڈD�&S��Lu�bXb���I��f�WdQٴ�jȈB�����u�e`�rT�Q�G���{t�Py�ԁO|�|\|�1L�#G�M��·����a��o��tF1�]�[rҕ:*c�s�%e�BK3=����R�.��t�y� �4ѝዟ���w�vsA*o���x~�)�T���E,�7W_q6�/���fL��o�)�����?>%b���^%�Z*<��[���C��Jv�T\:x��� ��5p�r\)al� ��~\����旮BNs
����ނ[~��%���tڬ�H�ط{��<��B�<���Ĺg��K�;��M����`����q�]���X�����e6ڞ%=�<͙�b[u�.���j���#{1��mL���ϟ�yg,�+~�X�;};�g�>,�;s�̔����q�����{�v�Cb`0q��~ڱ�����3bY��`a�`���_Ů�� S�є��	��F5�1-/�	L�e���"�����c����e\�n������
u9��9s.{����H���ŷv�Y�)+I��AB��Rk�q`��X7����v�J�8�#g
�$�m!#�N!�n G��L��*�E�8�I�*���+q�S޷�����W^~��u�M&�N����h��K�g����)�ԁ�:����x?��1�[�hF�Le+�[=>�Z&��	�fB�+wɔTꚪ��&!�F$�B����ؤ�^�6\fp�
X� �?,���5��:S���F�9u�qQX�i�QZ�����U`ڠ3��'�b@�n��V%Eqp�A��Tc*az\����ن���Ӏi���@���۱��\]u����ɡv�\�U6��*�Q:�|.�����g)I��Z�ό�J�&b�e��Xͩ<W)�t�e�b�Y���wݪ�t5v��H�������:-�GVZ7o�R-�u��wS�S�8.M��k�X��n�u�Y���j���P ��~�!���[��hi7B|��n���QBU�V�v��Z1��� B�A�Z1�����b�8�K<$0��>P }n�}d=��ʣΡJ�>J�=����Jw�:�������QS�r�Y�TV�=� (�@�Z#T��q��
�����.�Sc�)Z91�3�p�m{�)T�|aj��
��Q�E��l�9��̔���#��YtS3g7��'eZ�a����ܹ��P�Qv��عo [����;�c��=�{`�r���2��3	l����$c+G8D *��vNרҸ����-��R��2��/>9
N]�ڡ�z�k����>r�6���~�	�ȸdZF��m���d�.+*�������M��d��ֆ0�8�'�s��.OU�P�j�d2BG:��sgbɂ�X46V.]�)�R�Me|}����4�J��	�!������f�{'ֽ�Ͽ���@��nP�P|��<[ر���RT�Ch��9�`Ei�
L�W�"x���_��@���n�s�u;V�_�sH���A�7�����:�"��{�;�%���p}�2N?n���,��%�h�L��L	[紉���0{a
���z�
e�:����z�|4PkQ`��J��������(0_#o'��=
^��~/Y;�v�l���m�D�c�Rӭ��iJMc�Gs*{�A���dݳ�3�͟5���09]�D��u�9"0��B,�A3T�����鵔֚j�cJW^L�POϐp:�(;��v�`�I`��יI
0m0`�s����Zlrĵ�$����'�F���ϤZG���B��	��2�?[�L�� ��hPY��ɸ�J�z	�� .\u�r���r�wI?�V�w�8��[�o^�B��9S�����Å�-COJ��p��o{7�r��!N�h�o��D�\�C�I�;��Q�Q�����iR��_���r謌 �Q �сD<%��j��h�.�G��W�� F0L�7��q�����K2\,��,���fNJ��Y�Xv��=s*R�
�2�l���l�����݃�G���i�P(���`��F�?�D8։v8�P\?�����5T��+9�j�C����b|�+W��������W���GQ���?.�ä�%��V-"�
aΌn\v����30cRN-.��p�qǃ/`�q��h�H�H�ؚ�ZP6�no���ʁ$�b*���q"��H�^��ތ�m�Ǘ?���\�dXF3��P >_��l����Cϼ�~z+^{}+��&L��)'��Ǯ�G��iGҨ�L+�G��6��j�4F籄Z��n�� t��.���@�\ �y|ꃫ��+V��cҖ����� ��G��ݍ�{&.8�,d�kMl�s{'`Zg\�U�C��%n0��ҷyݶ�������2ˈ&C�U�F�y�!�8�DDt�LpI7)�1<p ��(zE|�>��N[�8;�^~�����x�wP��Η���q��$��9;��Y�^|8>���aͩ�z,,�a��B����[B�݋z(%�c�q��:�E`$C��ò!�(��әp��ʰ&�;�Ң�$0UA�R>%���'���D�hr<��0Jc�W���M�A�sH��#(��8&�1�2���eZ-U�%�c:�C�2��K�$�Ee�I�R�@�#vL+f~D*�����ó����B�fZ	v	�^ҥѪ�T��T�KQC��/�9�N@�7�̀�$�ɰl�1:'���-<�4x��G`(�$żO"m#�
��nY��A>�z��&�e/E��+`�>�(�.q�s
�F�uT_}%���\ܑ=z�s>�>�I�����u��駀J�V��sZQ<�wF|8m=,��KW���L֝�\K�S��~Vj&WL*U4�5TǇ�r?N^:_��y8~I/�1+p�k�xJ�\�8��=���y�0ڱa��A�S�>цY��h�A�� 0j�i��N�=��0����j`	}�i��'WP���9�g��qc ������=�K���z&��c�U�(���\*\Ì�4V����D,8bz��{����4Y �ݏ�r���gc����e6l|�v� zp8/4�v�i2#xғA�/��7��I�n�yQ���R�5`� �:2��x���Օ������7K�-^X"l��\Ÿ�h�r�[1��D�Զ�d�s]r�tQH������]Q�F�$oZ����F�Y��M��yt��ӭ�9{�4�z%4�B��HE����X�p.N<v)�/���	Φ�T.�3d/F�	A�����;�xi�V��ї��o�z�4g>�A��P�Q�b�ᦿ�6��#6S4n���o\AA�$�6u�x���`�;�s7�W݀�����_�8l�TQ�s�U��n��]G�9���^�|�]�"�:ґ2�Y8�\q�9�W��ϒ?���?cӦ�5���?���w`��@<�%�Jw��k��:��ٗ�&��bP��7�S��Uﬔ��SC���XD񶶚#i�Scc��?������vȕ��:��kAƏ>��v�����ە��8�=�����ODdʴKuu"�q1Ѱ�����J�@���b�EӢ���7�_�J!�ө�T�2�Xu��1�ʤ��T��)��A�G,�H.-sLC1�8�2l��ca��5+5T�ԫ�i"� J*��V%��S����2)��P�"T^ӋN?_����ҕ����
�rϳ��}Oax���S��K��}�.AwR���:~r�=�����,71g�lt�2�>Z*�Q(P*q�R]��X5�����@y�V�R��X
�KҒ��w�
Z��u��]�'2���V�2�&��K�	\z�J�{�V_���>��a;��Py�<r�62�
�^8'�+�^�l*���<��ۅ��v�X�"�La������Ů�Q���v��c�A���Zi�L������O*��Z�
��*EF�%i9�ԅ��W�A����߷?���t��-ttta����p��^�~#��Gwg����8�������[�� �ٰ_����~��J#�xf��R�eEit	.D�F�<��0�[ t�	�!ю�߅�]�1�'����8��eHE	Ly�i�^ZKĹ؋M������ԉSЙ���� z{:�|�"�;|2�]rfL�x�cl�A��{��JL@�T*���,րI�d��Z�hܔLt*�1DQAg��k.;�\�Z:�\b�rO<�<�����-[�)S:es��y`3�OF/i�A��h0x����mE|�g��}U�rP�M&���� ژ��.���'�R����~DPF64���竰��#�0׸M4b��x��7�p
�LS�LB$Jq�R'�9PX�hˏ�����S�]���II
�k(�B����g�=�b��V�4�);3�`U��EV�4�wN��Ea�3��hN�1�*�G���������<`*��Tg�RcZ�͏:���A�<P��B���	͏����U�ɮ��+�Q�@�P�X6�H�#L�옶��+1K"�:-&GM阪;�m�*`��, Luԃ�4��8��;`������ɡ� O��6���[��,��	��+��� �^qF͞�5j6���R�眶���CG�2j�G���F˶�-[.H}
 ����G��bRs5-������.y�%���΅O��L��!���e����Gu(�f�h�MՌH�;�]9�Tj�{����J����X>"���k��p���۫3�{g}o��;���_ށ|#�F�B��q�'%�� ~���J���_�p9��4`*+��<7�G��?CB���]�-����X*8y�;y�f%�WK��]��8h�^G��Z�R�d�ʨ��̞���]�W,��yS0��#�<�4m�WbU���[K/�E-}{�⺍x����?��b��,93F���k'M��ˀ#��n��>�������}gޢ�_ߩ�]g1{g��<4���v���y����u0��v(��XZ��7��P��_G)��kYB�ػ��Ł $�#Yo�0�л8 +�C�%zG�O��Y�T�j�Q��V�$t_v�B͊�GΝ�c�.��',ǼçaBw	sT�܄�RA9�^�����P���oģO����o���K#��@3�DQ�H��?i��a/�[��h��c$�SYDv�L�������||�`��Sr��	Y�и��C'��߭."Cۏn_J���2����� �Ƒj�c��.|�sy�Ȓ�)?�n]�b"
`� ��۞��\�Hj"Hʘ{)��J��E~���w��-��bbC�\h�[l�Q 5�'��D+�2�;�T��¨Sİ���� ����cUg��-[��@�m�z�sn���s��Qk�d~h���LRF#��>�֎3�c����Յ*�-1�p ��i�Py�O�A�j�Gd�u�c�˙_0`*S2qh�(T�"	N���g4/2`*� *5T	L+e��O# �ڄaA���SD��;�6����dQT��p���k����(���V�t�����1!��.>�&t����'7�w�� ��N�u��F����j(�	Jk����0�qF�r	��bu3��4^1P��#�2^X�[��C�F���B�!����x-���%�k$    IDAT^���q�=xy���GO����i8��8��%X<o�̵$u�����-��5*~�f9{����<��3F�D+xw�Jӑ.�(#-3��R-P*��Y<��+g�{_��e	t��+�������?���X�+�a֜�- 7����k�.���c����ZQ�g��� �i�	����(�Pk 6@ɿf�r&d� %� 	�fBy�hH���U;�|�NSB#�����������3���W��O:��qT2�t�ſ�ڇB2'��o}��I|�+�l�"���æM��}�N�v�q���c� &�"�!��ޱ�����pL���óu$s��8�P�2M3ʈ6�H�F��+N�՗���������y��N�M}Cx��71c�L,�5��ұ:R!u�؏�Tr�ɟ^9����O�;�̋�Gt�e5��%pN��J��?	���\(�Ss�QD&2�o��Ux��sE���q� �t���Jwaթ'����L9�/��6�m��څ7�ڄv�k���g�S�G<�3��ᡗ���_އ}C�+&��e�`V��Ҏ U����t�l��c<��٢Ԙ�N��H�M�PRҚ�1��ՋG��A9��)�b(�gE�u���Prh&��J�eǴ^�I7e���v\M�%S��s�&���aE=�&l,���@���0�;
.Iո�]��d��t�&N�*�[
t��$��ô�|M��?�c�9����z��a��kN��CR�S���P�����hA�Oo$(M��_~�\3�:D~U\�r�I��h���zA��h���Ep�_5�?sI���<ΰ�K��\C@�%5NX+1�uN�1�F H��f0��t0?:���{���������������vkQ��]��P��m|����~ϭ�.�RUf5Or�M���h2e������#l�A��%Q������>C5���<u�0{53C��5���/�鍲mse�۬VЮ��G�ZB9?�Pm�M�E3q��X}�
6#��Q{^b,̘j�<�:.I��,��<���lz{7^ߴ[����H��:��Puɬ�iF<� R���9�	����kz���=q�zG%�'�u��;)@�/�9����\��K7��xn��65�w�P
�N�'�Uc�|͈Eb��	�~s�{w�[6�v��[�UZ�@ �u���gN������c��V������R�Qѻҫ��+���KFY%?�F��p���LK��٧��������M@gHǕ	�F��fv�D��j@�fV\#y��9�g^z/o܎w��b�z*g�Ik��`�V]o�Sej�=� j1B�
o���P����#�7��:_� �S}�~(DY[m�|L�e���^\�E����F��H��x��ٓ�����q�	11稔���̜z80��'���c�H�t������T�x�W�]H���	��x��`�+^���+��B���JL]gV�tv����1�zC��G�M��Y�4T}�)���v��qs�5f�D;���8���4*������M6�k*yV���J�e.0^@��"i�,���4�өR��Ҫ��#>M��k�v�"�46��k�T
�ɸ�1彖1UF�O%�����+83��#�T`JS^��J`쀩�e5}��`����f���xy8k�����To�����7�$[h���g���{�Aߞ��֓�G�޷�ht%t�ƞ�2~|�x���p�Q�������I�`��\w�%��C�����j�h%��v�/྇����

���*�*�'��׿�9�s����!��]5�/o��m~|�=	\�U������^�9���O�wͼ'��z�����݅r3�:�Z�YO
�� {�8s����߫�J�1�
�8��.��������\׳���}�ϗ0�twE�z(���'e�^��̙�P���)P��x�nj�xe�^l?P[�}�8��Z���u�y����$�Xɻ��n#J�,f7혆����*������ǿ~',�.�6	 ��L��=�;������u�=9�Y�����Խ��5�W�[v�FZ,����|ud���uRF6��[5�.��Hh�-��e�\�����E' +&K��}s}���U�ѵo���E�����&u����q��EXu�2�$�*(�����OlA�͹�i�1�!]ut(�\#����u\L�YBg����%����H�F-���5�u�"��ĢG`��jA�2+�y��ه�p?�Z0G͟-���l�
�MU|����q��L#Q-\����똪7��1��Q�%XS�(Ӧj�n"�J	�kN+�����ء(�X�ٵ,����ۅ��n��łF]��JM�"�9%�&�khJ�1�dvӘ&������ڟ�P��̪�L��c:*]�D;��GbV�'�J�j#Ί�7�Ai��u�$Y3*�����Ӛ�C��W���!���{�2 ��X��\K,ґz�{�H���C�k&�$X�kG�Q\xQ�O��bMZ�7�ͷ��?��9\�����KhM_Jj��eՀ ���1�}p�S�hH;�grh���s�UV�Gr]I-h���eN_�Wnɚ=����4 {n�^"���^�p�xH=�F��V��8�Ny ����5<'�#�RҠTj��R��^{���~�0^ڸ�g��S��CRG���b�����k�4�s�[���՜��	&�ػ.�0>���y ���q�\��&�lL�$vy�%V2D�9,�J�R��fyTЕ
ᘣ�������ˎ��IqtГͮ�O@��3����q^?�,�7���i�<��Ml�~�
(UY��!�lRo)%�S_���2*˯�x�ӚTf����P`�%�^r��A9��u>Y@xS��_ ����)6�1�&#_O��<i@�:��)�Tt4���+@�9<҂��uh�B�g��z�e�g�L{����Ӫ�s�C\T�{);y��8��VEi|T:�j�z	�X3'w��3q��Xu�rL��B��I�²E]���\�]f��/
�����־�}���h�rhG��$F���ٕ��-�v�T
����w�t���F�k�YW3Pۓgd�be����q�G[}g��G��>�UM���Ε3���r�tHce1��G�<�pefv���yg,�Q����HG 1n���;�����"�4ZѬ�c윊����lg8�1Ϗ�b�p�|��{����_�w�j�Ro���4������1Gk�y�uה��r������C�C�Y�"�cI�4����<����k(�`�"�ۃh��T�z���!MH`�h��V�E��q�,��L ҥS�1%��z\��v��sn�M ՘�ٵ�^��;32��׆�����4?bt�Q%�q�RRS�DJ�>�Ɉx��
�M��l*���I���1�c��իU�/��5��?S�~��ݱ���>�|~q�2Vcrg��L���eL�K�_�O�;<���8��c���vWMu �ΔC` ��cy�_�z����k�?��h��b��h��\���}����9���q1}e|�;�Æ�{�bY�a�$���\}�1���F�?k�Q;j�<�nT����g_/�?��#��b�L�7=�5���$e$8:g�0J�<
EάŌ�������8[���o�.N�:�ZŮ�px�W1k�L��Ti2�*���v��RR_|-�o��WЊu�C%1KX�����>HX�`u�:�l�vC�a�ݹ��8�������SX��[;�mg��Ϟ�n� PA/l<����{ڑ��d��\'} ԯj�Y����g�ЭC<3	�6��D{�$r|�FĂ��n�a�
JkՋ��m�s=��Y*fS.��L)>,7[�)�`���o�o�����:>�8�)p֩��뿈���
aÎ*�{�xi����t�"���+3zѤ֒5��9�R��z��t��\��]t�|�rq)��lC�/`'�7H�Ne�=&���\?2����K���0X9. ��7V��[���hG3��rR�$xv ���
���pf
�xtp�}�k��g�%�F�iN:�ƬѪ�v�*���Z�$���J Z��t"3�a{��S�R�0��昆�u4�%q���i��άRy�:^��e��y]��6WG�F\!0EI�1�3����y�%���R��>DMS`�4�~�wM�aܮ�똧���3;sZYժ<?� �t,�T��C�4��hh�	���$Vb�|]G�X����we�j��|�,π�^� ?FKT�-��]Cv\�*`_tV��9$y�y{VCW:6�IVS��11fq3F�3��:���<v�����~�R;ݯg(㰧Rp�u�w����^�VE�R�K�@��:����7*���pz
_���X� +�)�9-0�,�R�������.��7��ώb��H����P�;I�e� ��9
�g�e����y������j tX�z$�b�/��F|wE�k���6UM���C�Iz�VE�R�!���h��Бh����cq��#1kj��;�w�8�œ~��)��:8�NX^&��o�H0��M4�G�����Pם�o�t��G���Z��E��-����uOk8�Ad���4Y���\���([{'&�"C�$�ua\�Gⵌ	2�r��a�y����km�:�H�\���{�w�ՉA3�#� a���ny 8��t]4sNW���z�-:�6Jd�0&��h�Ց��7'�X�3V��GN@�5C�$
�F�E	e^8�������c�x�0�B�.���"40d�6�h"�h<&�Z_OA)�<<Ӝ�����E���iY��ێ�����t���+���E+�y�TƱ��򻟱A�i*����-4���Z��iǀ�(���篹�;k:��^2 ���wg���q����JOA8ՉZ;,S�W<�m�Yȳ��ckύ��"��QRP������-oF��5�K!]�`hcqP�I0z�o���-)��(R��4r��m�CF߸�h���l4Ћ�3�'N@�&�a�1e��Jv"��4A��`Zˣ������1�pW�\y���S��	LSqdYȮ�060�z���
�zH&���iMFB�3���1��C̏ꥲ�8�/O"�N����l��Z^��t��$��3l
4�B�V'�w:���GO�T���a ,iN�:��-�O/��/~���؉�=q|����3V�#��ʝ����SO<�5�O��|���0���$"�9��b��w��`�6p��i!�(��/�?��ܲ�<�w/g�>�����*�ň�`����X���E,	FcbbD��DA)�P���3��S���>����w�OYk�������g8e��z��}�������:\w��9���\���L������?�׽z�h7�l^��q� S>�Zu
�-/�S{'��֣0��Ia5vf�3!�r�]>�F�tl l�e@[�𙋿���<Z���O���l�T�.$Z73e��1��V��j��쓏�'>x.��-+R0��&���0�q&��-M\{�]8��p��(���
jr��4��3;�/�j<�#@�)�N�H�
��"��>�Y�<:�]�\��˦�R5]���9�G����p�ACR5`��ϫn�]�>��]��;�=*�C���SU<������`�0A���(&��7W�?><�����eg#�ŞZ�t���*�5Y��J���:��l��?�)x�AE�/���FUH�\,�vu��-�g#�U��m��5{�^���?��+*8x�oY?��~�O���M�I:��� F�Z2L>��� ��F�.zm����
f��C��3v>�^
���t���I�:�61�e�c�m8/�!JV��+�=`��ꆧq�GQKXhtQ�C"�m��4��D��|	>q֘�;%=�R1,�l+Qn!f`�?3?ʈ���ƌ�0ŕwp�Jyt3��!�=4���	Ͷ8��.�Li&��Aq~�"Z�N�}\�i��
���xYQ��6��b��
0�s=��5��I7���>)��j� ��ݕO��KkL��j�/2̰�'�/s�J�&�ψ	�#֌�>Ivм�&
�r�\=J�i1|F�e$��DUKq������7�`v� �
�&\���,QyI�%��5���Z�d5ћ*�Bb���ҫ)�{��g}3�\r� �M��.ERO�^�V�}-]�4�ҧ��-2j���I�6y4\�
I�1Ɛ����ؽ�����8��,8�+���}DU L�����/��<1�03�n��T� ���9��S4K���Ӂ��$Ц��]���.�����<N8&y� <��vo�)��22*����c#3�����'�7<��㘢 ac鰆�RG�o?�����EAC�ML7�j��v(��J�nfشy+x�I���&lzz+m�2��A��e���BGAp�\."�4~��!�`*F*>W1if%�zo�]a��L=�,�����j�	�zlY�+"Db�J������o%+�^jϒ\��ס����=K��8��)]w�X��Rg#mX����(�Kdw9f�N�/jߣ��u?v�5A)3s�>Zb���n�.ഽ0-�hl0�SO>'��(z ',�c��y�6�_}/h��(#��gb�K�����w>�&f�h��ȗ���L6�F�\0�$�rKVڝ��%�l��ɧ��*1�%B2�	n~}~^A'X���t�E�>�M�ܧE���(�ש�W�V��.�ͺ�0�r�[����<>��o��ox�ʐ�V�$ќT�k������W����,��A]��T�Ѹ�rT�>�3�:!��87��,�I���g��+>����&%�Xn�-US=����	7�R�h�s�L4͠��i����r�z�C,"dD�D�so6yy�"A*���� S��! dߨ������jNVL�a�j�Z]��vgœ�	������,��J�i��S���i������)n7����ĕ�ß���qs`JW^i*	:�b Y�>V*��"#�<g�B�l��s��Z�5�����3A���{�k�������0���T�����7a˶��ky~כ�ӎ���s�f�����7�ÛN}���>�Ib_��2]��"�<������r_�Q�"35���Onŵ7>��;[�_�m��Gz����Y�,�����/��UX�؋"�Z�������\x��0@�΄��t��a���$a��~��8�ͧc�q����|�ﾋ3y4�����qIY{i`�r���kI����w�^k{,)�-��sN}V.� oU&�_���s�M�݇�o�I�=o|݁b�O�H�#���S���jm`���׾���2�T��/��S6���<�=�#lc�B}~,�k�B��A��p�����o?����|��݌��|�}a+��.:�l�~�1�})M$�{��տ�g��:�9do�]V,@�S��A�>&f��/�[�;��dd9n�x8�#���9�X�
�I-{���Bq��8�C��d��s��'�S�w���}��r�&T}��S��G��_ߌ[gtb]��C�Ʒ���8p�1INi�tビ�����m���ٔ�y�,G���+��nz��t�M����ĭ>��J��T���#�ۘ��I<HþV������O�����QG��8�W�?���{��S�ZH���n��gg�+���꨹��C�^hݠ�l\����̥$fFlH��kK�0 �YsI��hwI5����VLh̪��I�����Q�V�F����'U��f�^��:Zt�e���0(�E1��J�k_@/o����X2�4���G{�j�br�q�&�~T�W�df���9�����W?-�E}�/vN�����	a��BQ�g_0I1����21�c��Y����cj��f��ѩ5ѧ�TW+s����.If�PD�͘�E�wK�$������U���7q#��0`*�ϕ�6�G�W�0���� U*���� r-��tЬ�[Q��,g�\�5�w�$Ks�&�q�����Ɗ���'KS$�����Q��ux��	t��e��sCS
M�N:4    IDATm����$�ߊ�A�#%�U�<���ŕ9|8��f_���}	�#՛���Ί��d&�����j}:2F�D���j�#lא�6Q�t��&w��^}�~X�<'�F�ˍ�0v��but�l��ێ��yw��0&fh�@�4�\a ��Y�ih�VI��sR�i��ɪ�L��������M���(^�v'�(�oϮ�T��*Y}��6�x���=�+N�b�Fɷ��¢�T�,#zb��K�^�@�<S��:�d��o�j�<�*��JCN���6OWH�D��\�}���T���{�|U���$|F��p�*1K	!!�@z�8���9�&J�V�6��N8'�p8�oV����WI>#�La�!>;KF3D5IZ��Gp�Oc�tm�p=��bVZ��j�M)���I�z�WD*s�⹓�>�ڞ�n5U�ρ�L?��t�ѥ���dN$�W{(�!��1]��ij�E�P��N��!�_Cب�8��~��3�3��nC�7]($�}��)L7�_]�~y���1O�Z���Ft����f֖�
���"�����{%�s�˘�A�}�_���c��뛋�H����1=Ѹ]���8 E�Z§{H$��ǕS��k�P���:��X2�L��sL�]�d� [� ���P��Bp�)�	J�+̧R."3:�^Au�,��Ms�~�LsH�ۘ�9��R^��d�)#)/���eԌ�D�E�9�C縘@�i�%~A�|	���� m[���T��J	�VL�Ń+(�L�:МG�=���=	�x�밬��VL{}�
���㊛��ko��|��ş^p� �J^���[g��7߸V*��\�Y�ZP�I�ddQo����E'�+$@�洏��I�{?�W��^l��D�E�A�L�-���_��<xX6+��l��K���l��榷c��
��_\�����3ii�\���v)�p�m�/4�j�0��Ͼ��_�<�>t_��)<������DC�r4#�q6�"dl,=�d�r�!gX�6���1����Wc��qiT.p�-�M��Zxv��%��
��;*,��R(�M�ب^� ������ϣSE7[@#��H�1�S*t�kz���O��;m�C+g�(�v�.�q�~{b�\�B��'�����Po�V���ce�9`O��nX2�TdV7޴���^�;��X�t�c#ҟ��>Wmc��x��s��N���r(a�("w��R����UeF��i�Z��Dv������w��h���G77���3uv( ������k-���������=�z� ����o�
�yɧp�!��,�+v�#u���;��fh?,��#t��ӝn�,�d�$�B��J��-u�9d�5,��G���˗�bph@X�f�: �*���9\s��xp��jwԡ8�5Gatl@g.f�h��/4Pku15��Û^��OmG�[@i`TgYq�	�o�4Ɔk����y�GEKFen��y�<�Xz�T��'�f1ɳ�ZT9/��T���Rޙ94�r���ap76~�%Ⱥ����W�s�����ZCX��Yo"�/��@y鈰x�3f�o"$hUk����1%0�7+r?0��Ԓ��Z!!��y���n�	@%�ɪ��G���+ RY ;i�Z\�*�!�^)�#M���N��(�Qj�"=�v�9��^s&�� ].��fH1A%	�%�NLD�r���$�<DOvREw,�dBûJfU�W�5�6gR��W��e�,�˲I�cE��E��w<�N��[U\@�����B^�$����
�o�����K�c���d��_��T�q�8FX�7	�'�t�k�.�����:�!�*�RJwK�-R��~��$b�-��ݝy]�'�J��JO����U=�Ǫ���+��H"��eU?M���b@ (A� 3���(1�KuѪM#hLa������7�z<�;r��"�:eF��P��%�T�l�⾇6���cOo������ӽ8W� �qhR��H��G���AgꚔd�+���i�D+x&��ұ[k������{�P�8��Ǧ*�W}�*�M�6yZ��R2	���K��ㇾ�w���v�y�VҒ���_ח��b�פ��Zm����Sr*�$���O�y���y׊�+�"3c�<LU�h���+�! �D&���	P��B�:�Nc�T�Fr�{�1u�x��'`͚�18���Ȋ�4����B����qs��p��ԉj�~�">�B�|���/�[ɇU�p�QH��z6���jyV9_?�<q��H�I2Û�>�-;U֨yP���\�m�g������?��*ОŪ�,��'��C�:Er}�*�G-T��S�`�<�ŏ��UzN�Y��"�|K�	.b��O�y����1�9�#N�{�z�~���(�%��;$KlL\����QC~�����~����f��Ez�I�p��D�^oZd�r�bb(�bh8��+����b:@u+��Z1�Ŋi��ԥ��s�|G����0P̣��s���Ղ��Gԥ�LymB��
��4Owr�w����m� �b����Z,��8�E�7����zDS4�����^��Ť���x�
��~)<3�ǥ?����n�[-�r|כq�)��u�̖i|���u���SN����g0X���E�+�Mљ�\�ɍ�k���P��G��W^sv�l	0�7k�g	LS��߾�C����d��J<�!�����|����5(I�Ka�i|���nA�E�ʦ14T��k�W����K�������<���V� 3 9��+y.g��.l4�u��U���y��p�fPZ�9��}K�L����>���'	�B�fEPng����`ΪC�#�~��%ȍ.E�ɡT�D�����f�ZQR'^��{�;����jU�"���X�K��c�Q���M�9���A!�C�M���.�����D)A� $_�ݡ\��݀Th�d�UȲ��.Z\�6�G��W �w��:�B�j��9�{��{�j�q�Xs�>�������
;'w�s>�Cpƙ�cŪU2d��g&p��`z�*LQ�0��J����ԓS5������ub��E��E�XD&�gAC Lz�i�-s43��G���d�x�YC_ۖ���~��r�"���fh��39:�fTk-�G#����X�t�,{5��k�=Q���j��-U04����Ҍ�ʁ�Os�TG6�R1	{�0��Jw����W�R���q��+Si�� SZ������ɸ��e��T/�b��G�V y8�yM�Z:���W��ry����S*�2r�KV���Z �I�#pk��B?#�G����Ty��-y��V.�UC7c�C-N.NF^R֖�sj�d���=�ĉ�Ғ5��y��Ss��R�#�DJ+���98i�%�"�5b��"�
e�L�մ��(���c�<�o2�I�%�0S�����$�49y�ᑬA��Ǝ�tr�ۡ�����5�:TΫ�
?[<���|롖oh�%�>ILH���U��5��<�{���n��������t�q�F�X8�>�w|b���&ܷq�ťi]G�-�e"���{�9�+~^c5��
^�J����Q�Ř�˹�����CY���}��9�&��۠���Qű����a ���f�^��Cv�;�r2NxվXƑ/�#/�V��I5{�9֪,��-/5���q�����[0]��2���0�ْkbR��Ϲ|�����Hw���>Inm��8Tۚ�d��SUa�y�r�	��A��"�Ԋ�0�u�'��b�����ئ���$K�����Z5jО��'�4��$DL��I&���x����9 UOo�I���穀Յ�N���("�Ly�$�6Nv�ɭj�b�'��/�.Wy6|V�G\��;��-L��pf;Щ�Lo�`�xұ8��Sq��at�/�y�c�[�V���LU�݆+~w;�~p��7��Ȕ8������$���K(Y�U�\�G��KX�&�S�Y�z�h�Ecd�e6���
������'�z��)��!���tK �riVP�ܮq�4�t񉏼r�1Xf�4:F�ACdP�����?~�*<�ia��4-�e&M鼑d�����*c����Gr��=&���lјeQ ��'os���YV4�Y]���]��%=�}�����
�'�p 6�@_˝xm���L����,]�^>/��-G:�NW��~O�i�q6���Sq�Ng_�JNY����,�i����I�hT)sLiZ��⇂Z%:��4���Jy��@& �,�X��,~��9���r�j��m7�
���fQ���N�_\p<��m;���j0}~
������7ߍZ���V��O��V�}�"%Պ������u����W����)M��=PP�v����8�e����<����gw㷿�!�m�9$���epٿ_�C���/R>���"�}dË���W��r�>��w��7�:����{z
��v'^ܺU��`�?�?�h��
��*��vq�����,����qe�����=󘞂��qv[��Y�Eka���M�Z-t�-��+�%"xٞ�l"��2�Pn"�]J�ʘ��*��t��㨌/70JR���Ā@���R\������&=��I���n��e�`�	�k���Yb���u�-t��;�h
J'�p��t�����G~�r�y�!�S2��E	��7�H��.��kiW]��3���� ���40TJ���
K��Fu�&UJ���*ccG:[D��G�I�~�z�4U7�z�8��/�����g'1Y��~��q�J%�K!��4��h6��r(�'Y��Z�{I�4�M���ڠ�_l�C����3�d�^����J�Thi0R��E'hh=�G�]d�(b`h#��RI���:W18D� �>�E*��_�Rt˙\��c�u`Wb%�%($�a�u��6k5�c#X:�t�Nڛ+�ʤ�\A\9��t+ЊiuAd�\;�%��ҥ��̤b�W>ͮz)Dӹ1?"X��tƀ[�X��W�I&Ӳ^+�
x��&�`O�DB��jL��b��J�0�"���
T�C�B#�y!&D��Өt�(n{���D��ǈarMJE&h$�:}�a��T���T��=5��N&�`;���	�'W�}秀�IF�b�D���+�Z,Is�YyL%)W�j�Ħ0�&H�% C!�># ��ţ4�PZGA���g4q�.�8i�r|�����p����>n��\u�]�:�B�F�*�x
�NU�e'^�1����( qɴ�B2� yN.�O�gbI��KK�X�$ll�%�z�"lK��RT����ǊgFb�մ[h��6f�`���q���{�q"V.S�.�����1).������=���&\�=x��1W�H�*W�$`9s�G�e��g�>?Vu��O��^�'�o�m��|���V����~�XکՕyWTm���JG�L�9I��@�;���Zd�L�Qk���'d��*��WIE[7����D�h{H��
4���}A�g��etJT)ս��螸�^�b��]�fj�"��ER]��"�E��(��q5�����U��om~b;���h���i���BG�7>p���#�����A�h�����Kp����+�b�S;0ߦ3� z�"JC#(i��M΢i�]���煙��|ڨ��r��-�.��sB����
ȜO!�������#c���~a��Vu���Uzx��N���y&�K�/��x�LS�2|�_���{�C/7,yۮ���+�~qȉ��L&ҧ� �N��guՃ~����L��	/��hē��	-�m1�S#W���m7�㩜�~���	Xws���DE�X}����)c�8ǔ�4+����.��v�Ug��N)�w7슟Fs~ArEʵ	L��"RìZ���ʞak��r!#�����4�ZS�)��L�Y#�S���U-���4�j44R��9�%�ӕW?�Uk��c�E��c>!>�$��<�9�b0������;��R�`bK�D�R�~�O��3�w~|-~{�X�ձ��K��}�9eL��,{L��s������W㒋?g�TR��1���>:�$C��kx���U� ��靸ꚻ05������f�X�4��]��_Yc~ӯ��o����2"�Q��@����x>��wb�Y*lʇv�9�*�b�0o������D�G�Z��[�����Jī9o0�%�t��i�h��f:�IH�,@�X��
(����.�J�er���]���.=�4҄���y�F���`h����HqV� D7HC�r>�MMh��r�N������:�=��Ö��a���Z
b�!�`'��)f��z��m�*������q�lx����=�d��(��!�cOH!m��4� ܓĈ�5_��^F�6��I�/�5��#�@L by����I3Ȕ�ȗ��ĳb�j�P���M��E�XDi` �.�hP^�V'�|y��q��.Ut�e��o�f��$��M��j#l���v��V�)rj�q��6{���ŻTQ(a�G�
(����Q,�D�X'��S�6l�eqp͔˨��J�%�bI�g��@���谄G\ެ�@�Iz�A�VL���2��"`�|�$G�<ܘ�3�7`Js��ʨ�+�BV�M��5&23� \XW^�)0Fi|D�-�┻ъ��{�!��^
��VL���]Me���]������3�kT�������4"J#GA�a�,cK(���:G�u��&����r���n�"#�̀���8n�}�"�%����8��[	9�<�� :�d��@�˵*[TP�X?O��3�|F�0h��g�&G)x�.>|=%t��lʵ{$A�=������ �G�����V�J:�*����*�g�7��f��F�H�׫c ���G�5����p� �Ï?�?>�8��/� S��>�z��m�CC�
)q���ʌYӹډ*-!BR�sp	�����$@�l��/iO��bՉ�dL�9 �	�ϻ��J��,�K�� ���- lLc���c���tN8zo,��n-^����ΚC��W�;�{�o�{d3&g�hu3B�Q��/U�:J��a��鍏�w&I'O���L��}��x�P��OsZH֕�E�����JfD㥢�KT��G��Zwb�$D�W�|޲�$|'O�u]8��׌��-�]�*���{1a$�i����Y��~����n�7�$D|$�}�Z��Q�2���~r0`�Aㄍ��^W���:OW�'<Rd��GQ����4����0�vc�,(�G�8�Ɠ��i�;
{,�I��|��c�Z����[�����������^@';���r�FF������� �룋�����mF\�8��4�>q�L���o����JVe��Ε7�`�l�ĪJVIMj,������A]��z�)�1��yoz->��7b��2
Aő�=����~��xj[�0]�����Q��0u��n���p0m+�
<N��4r�[���U�8^�ȣ{&�3��U�s�^�o���Q��8I׬�/�
⍭^�Q�Z�oZ�:6�w�*(ĕ��\�e����V��qB��o���0��2cm�A��@k~A����$�h\��G�gƘv���X+��0�܎	�¹�$������:w�b�$FE���Y��aZRQo#h6�f�O��,͏��4rI��C\��`'�^eӾ��v��ʝy|�������Mt�/*��>�����57�!���V-����v�s�a�x�<�u߾��妛q։��_��TScSrF���j`���AlLC�����ꏘ��:�B� �ib���w���}Kr�Ж��9����MW�^g�����uN>�p��!ޖWF:����|!x�cz����_�z��z@'��$?�J�V�lN�]�~�ڬ��s�~8��}0���S-�;�L��
�ÞNMX��`򂀍�ҿ��Di`6H��6��di�0��K�Y�`�s��d$z2�"��������4)w���5gq�^˱r�0��yi�&𡄲+�t��q�֍&�8��R]���Z��mv7���I�:�g����E
C�8<Xd���D�$��a]������q    IDAT�y,+c�%�rR=e���Zͺ����>,,T%l�$��#9SqH���r����&�Ah��Q4N�I�cj�� z�A��%]�<_��ܸx�2��-��fP������x�k3�ݬpi)'b��`�~Z>?���6���4���L�2D��\^��CH���4<&}�y:�$E+ɞ9+)�U��yō?���f�Ǟ^R&����2�Җ� ?@��do�\_L��+]&�@��D}fV\yyX��QYB����Ι|�!fY���Ҽ��L+@@PZ'0m!�ˣ42��؈��E�T�j:p���饐	��L����J���&*���`5�8��J06B�oM �rc��[����s�K�q�,���zh��`�]I��@G?YL@I���б���̄�Uc�{��E�,�zV��
0�[/�!�h��,�, ;rHJV�|�U ���L4��N�hn�)L��: _��a��rӵ�׬�0d�z�=���c�K�GN�k	p�F���� I2,7]������趫H����(��"����Ȕ��+�O��4�ɊZ|���rQZ^$w��"�Hⴌ>�U|�U9ݼ�,��A��r#��0�d��^	D٧��5��U���D���A�*Z5VI�QH���1�w�kq��Gc�n�A��=RU(a$�اr�d�_{/���^�	�K���/@�$��ue��.�F�Y��C�?/���^�������+!������w�����9�2�*�&�����DF7�*O$]OT�T^!�"ᬹ}�D%�*i�Ҍ_��2C<���ug\�Y���IB�wl�Q�2[7��N�d�VJ����R��k�ߑ(o{X����-���x8��w"J>m��n�DЬI�j/\���_���L�~�Q2ڎ)�O���A�[��T��?m�W݂�o} s-:��!UD�0�\�R֌��x����&S9#s'�1��`[c����pK���gP�k�x��5��Č���<��()�Ą�����}���<��]���W��:+2d$�ı��>0�o\�kLײ�f�K����P���6p�i��P�q3�~Ll߳Olf�NIM?����T
��'2ՋZ������N戈ҵja^�o�0�>a�/�j����覅$�J�R.�BAq|)�9�Z�I{sI%FS��v�Y�f��-J̵��}�������P��R�|�Ns/M�C~�ϣws��2RŜ�c���JD���3��G����pJ?:�ӕ���s=w�uD)/�����*�\a͏�H��Q
g�������h���W�A_���I����J\��N����8>~�;���R*���)|�R޵�ଓ��?^�7RM]L%M�S �V_��~'�����NL����F��F:�)��~�S^��M���7�¦��e�U�S��*�X6��I�Y����Tv��(Y�T�7��ɔ�4:x�y<��<�i6<��f���8�3��Vr�
��ĉ�{�Ь͢Y��펿��8d��|{rl�¿_�3��s�M����M� �-���B�v��O_��M�gË�4�j�VMv�뵤S��\�!-�iSǹg�����,�kVFٌ+to����_�k��,���OO��8�G?#�*����������[11ϡ�4��A0�>WV��8W��=�G�7�]x6�>�PC�ɖ�5u�����Yg��Xo&�GC	2N�<z�Ϸ�:*g�U�z�&���v�;���ȗ8�@�ssy�;4���O�1\��J>�	��������"��-��>:!�/�{�kʚ�/��m-W���3�f'��z�0�tiPdҔ{J�5��R2�!��.��5m���H�e�RO��D�N�cca�y ���0�6Z���n4��Y��̱O����^1�o:���]�$e���>����(����,���#�`��]9��)4�������7�ײ��h,ْj�&܏ڷ�I��ېb��0ѤAYSO.�$ e2)V�g��z}%HB'C���֛�5���S<tޓ����Hzy��kb�.��'��J�(�`MV�i�ӕ�If����C$��BQ�n�ë�[�g���D�G�1X��HN�?'�I��u�Ԑ����Iބ�6Q��;Z�u�@{�qW��#�.�Q7��8�n""�*���ba���^(J�n��L�%�?�J�Þ�B����FaMG1:���D���-YS	 �$�wHD	�-����~'�Ti��M�}����������:]�#)�j"+
	#����y���X����N<�x��8�1�$K>�X4ٿGPJ�Ӗ�B\��^�~��8QC�WD z6��;'�/Y�R�('j}�	��	�<�Ź�D��<�"�7�a!=��F��i/�{���e�^����i�\���2h���;�RM���ۏ1�����b�EY��L-9H�����'�Z��=�����K�Eݏ1���A.�� ����Y��N1��䝨�$H)Pq $1H���=
L�9�0[X�H,��j��X��BއV=2�(�fcͅI�=��\�y���8n͞���o�Yl�j���S���1m�cO��k���{��|PB7;����C9+�B��`^�w�'�h#K��C���%6@G�>�)A�&� �^���`�®����}|M��te��+�x��<4�K���5�b|�u���՛올b���x�ٝ�3[��8�)�X��I�<s���S�-�������?_�nITG���� ^|Dj���TϽN�O�N�F�>�Ln�Ӂ���I�T V?��g��狽v��c�<J�y:�+0m��d�lJii6J�ǁ~Z����au��8ߝr`�K��YR�HYkN��f>�J�(��Ĥ�Ժ%G`9P�|����*A��{@�)����6�Z2~�$!�m[[�Vo��'��,�)[���^��l����9�R8���7�#o{��0}���W���`���%���o9e�
�{��\���a��k�^�ϊ�W�z*�L��O`��靸���Bt{md�u�"'�}W��g���M����~��OMJE�јC)��1G�^�;p����`Ig�I�K�ؼu'���Nܷ��8��Ω a�����"�%�+����eZ�&0��u۷<�nc����O��U?�����*-� />��$-�c�}�F�B+g�'[�W��7��4j!HQ��Q�����O3�/V%�mt[�+���'ߋ�O\.�, �/=T��b�����' I��pY��X�+Y��[,�9b!z���ؼ�����h��R�٘��E
��>��R_����I_���;hr?�n�H@�M��b1Qg����{����:�s
��߽����l޺��f�n6��@A�t�|Q$m��Y�N���c9���#q���`��m4g�S�e���d�"l�@�6���}�կĒPs�A���{LI�<�t?�r�j=�/7�P��d�[���nR�����H���0J�p�rii�g�c�Ry�^���J��/�t�m��j�T>tQ"0&O�.o��W�3�+��B���c�`?<���9u����h�S4�i��I@kvAW������S�����0���],-���c�>	^ĺَTo�zU�����Ӝ���*D4'�,�X��D���	�)�)eֲ�tX�26_�*���G�x򡱥���DO( �D�	� n�.	�%��
�.�DB�=�4��(���K��g�����,�F�B*p���{�)�IG=k�}.	E��NT �Fq�IC�c�	�1���	��t���M�l`O?Ga�dV�J�M�,
P�2���y�*��"��.1�M�.e�L&$k�6KN�n����.vBVy�&�!-��A .De��n������)��p����o=�9z_���I#��L�,�Ȫg�?�����^�Mw���gw��љ��4{ˉj���[!V*p�ja"��zy���b /䉽Kk�dE2֛�@mD-��%����I:�?.���Z�x��t9�M�\+��R��ZeF?���Մ7�bÕB��cS��jO�i�mҽ�dڮ�#�D���H�l�L֬;���s�+'r�%��N��HPX~0��Q	��"z7� �&kĞ��g�Ӽ4��2��G�9��>��F�xۙ��'���]& �=���fi���d^dl�t�/�7��%�y�WDn`�l��Tt��19�R*q�׏����>��
%���/�$�D_��j<j'Y��5(^��W��#�WN�x�k�}DpE��62}V��gq*�r�<*� �@O|/��Lo�y,\�8�(��s4)�եj�����~Lm�0�s�׾�di>���*���5�Ƥ��,l�{���|,����\x���y3���9%l%6�h2��N֦ɢe��o]�07�2�������-V!���d����G)��:�5��2?���Q#��6.F]�c)�8��/�Pa+W��y��6�a�X� O�1��W�)?���0M���9+�����b@UV� ���w;=>�8��)�"�$(�1�rw�x����GaԌ��K)/A�S;����&���^�?��x�I�IUԁ�e��9n�y-�|�q	`���1SKQ�k���Ky�T�Gw���݋ɝV1�Й��U+����`�Uݠ=��<Q�.�5jBG����:���1�f�J���7���vw?����7��''Pk�b�!�e�ryq5u`����T�0ܼ�<��՗��ߌ�?{>FI����g[N���\҅�ˏ���P�V�<��BU���6��?��ܺ�mJL�P�U��Ai$�g
]J��{�5����_�8b��l�.#���5�MUbQ7��_��mW�7��i�[}��-�/�]����E�8� ���4����a٨�C*����s��/k(FC��8�t 1�� ,�9�3�9ޟ� s�aݏon�;��6�a�NV�:|�%�n;!�v��Ԏ�8���ԟ�ǿj%��k�]{i	f�%�|"'���.v�ہ�a�7���Tп��=3�n��f�+r��jg])ZaI�09��DR$��d�*%���etēcH�`Szy
0m�. l�e�H�<2$=�:�U͏$�a�lS�8s�	����A�l����J���,�^1+v�乬��M���A�/��D�|�������$��u�Խ*,�WYw�dnj��!f|��U�K��g��ʪIh|��Q&�1�J~���-r!�UGl|L��T/���Hk_�ػGɍ1��c��)�!@彖�^ca�\JGߢ��>�Co���GT���>{�*�q���,2�2y��:�bh$9�����Xݎ�s��X��(2�I��&�'���Q@�|�>�9�J��q�% �$V�Q:���U"Cq��U�=�
*4���1M&5��������D!m=�J��ŖY�i�����>iqeoʘ���v�ڳ8l��8���q�IGa�=Kü/I~-�#d#�3}�v�c�����3���hv��f(�ω���[϶$��h2K�/tڿm�9r��a	�b�����D�cb�.R0,�Ǿ�cU�<����6:E")���>��z�u��L*90�g���y�Z��%}����p,_V�6#�%���	�F�3��5Շ��J�Y����OD9%Z8D�[�|:�S��I"�+׎�\��9�z�	�q(v��12��(S6h��NHi�j����hc��
N:�P�u�18�1�w����ϧU)}$ []�-��ww�w<���~~)�0�%G���%�r�&?�W�LJ� Y�1x��U���ټ�9y� )����,��j�!.�u`����oT��T�E�N�6̹� �k�PՐɕ���#l�̵hQM�D��m�e��<n]]!�O�k�V�GR�)�y� э>&��1E��=I����\W��ޓ��A��l�5';�ԩ^����6Am��b	�%��4�R^~&���T�5U�e�,aW�]��`{�(���@���J4ǔ�Z�E��J`Z�a�Rް���ItjL�-��Qn�U�\�˜KT��㑰'F j}90��S�F`�DP�ǚJ¥mʈ��aG`�
n�6�J�|�9���#��G@�L�����O����?����M80=���H�)��3[f��������gQ�$;�=�#Շ�5�BwM�^Ό<x��*u�o`:3�Eu�UL�ܳ����ϞR�A�ϊ�.��+�i�,�N��e�i��7�c�����L,�� _��_w�F���7�mut����%)#8�#�#>1���)��\��)<��c��C���w�q;:J����$Y�82Y`�;�O� &�vZ+��TZ�����e�yW��0fZԄ3�d�wR$�LB�*ҦP����س�/�c8`��̞s0�R���� �S���$"�I|�(�M&�1��g�i��_݉u�</���\�b^����i�"���=���?}��A�FTQo��j��Z6���(��ŕ~�Ώ���I��쇧�����Ãvb���^��� 
)���х���0�<�x�A��gޏ�J!��U���Ec݁<R���_�1b�KX&��pp�G�gl�����q�#[f���tN����Cs��Qd`&���~�[�J�4���<B�21
��4"�eУ����Li ŀ�(�2FK~�� .q<0�ų��$!	L۵*�v�BY*�e�t��a��.��-����Q��<�9�����F}Q�Jx����e����^�uu��q��#�𑣴�JMV�b�R^0�ɬ>s�_J�n1;�@�,u�9"��}�ł�L����՘X�԰�V �,o��]�Î�|i��X��B)e!�#&�+K�פ9�ݳ�M����E}��QeX~��arC�4:�������9�^�Аjz���M#��.D�KvL�=��[��<F�����ƍ�lC�z�|�gM+��,N��*f�1�"�f̣d�!qv2���Kd�#���QY<�?)���K*���'I?�5������2�*�M#.`��<N{����cp��`K��wx�'��w���S�t�7�� �xn��#*hw���l�c�H��T�$2j5���d3����Vy��;]�J����
t�J�����k��˽��U�LV$�Nj�q������[_��J��Alf�N���
��_IrJ�1^O�L��JV��8�_�>�U�l�&��OVJ)q�G䅵'���ħ	�R�{�B����p��.����d�����_��m'A�Ұ�-���
��RÅ+�4q�e�AK ��h��ɟ-6�(����A����p��Ǌ��TX!��1$FH+��ҧ�}�.��x��HGQ^&c��9��)���C)*0\!d���Z�DZe���"%!e�&���x�ʜ]=F�y�g�V"mIB���K�O�-��qT�];�G�BT$ޠ&GdlE��	���y���_KM5�p�9��`���.U��X��/��+���]JKr���4c僁Ө��[���e�ZİV�]b�dY�x���<�zw=��O���u���_{h3�#0eW}
f�����3�;��B*�L�u���vi�Y)4?*�p枔V	�uS�g#`�R^S5?*V�.�u\�l��/kg`�5H��VK�y�T����9s�+�6���'��+��q1-��
0���S8�s$�|��+<p�L�����w~|���nԚM�z�����CP�j����s"�]{Í8�����:�üH���y�ei�+��$0����p͵�bn��F�R���V�.��˾��W�D#O܇6���]%�L8��,V�g������~�H�E�h��)�eSY��l�����k��� ��R���,w���
�m�쭐I�>��?������{��%_��8��3>[q�ѐ�bѐ�R�^����e"�i��%�����x�g�	0�[*0�^�W�{��� _*�P��:4ꂡ\���~��b*Dga;�w�������,�b��P��\����L
e�2a���1م`�!�=lf��3��n�|����;�B���� Ɩ��R�0�Cc~a��&p�����K����_�M��
f�V���&�?sqo�t����TF�}���i��^O��MϷ���C�0��{���nK14\A�VGmf
�S[�jM��7��~�B콇2����&�����БT��jH�    IDAT�9�"��j���`���܍��~a��^��0*��=�!�[�OI�x8;��"��! ��͠HiH1� �M�q��=*�4�+}���v���
�2�F�Ӟ&�")��x�uڗS�ˊ)��Pʛ-�10:��Ȉ���7��4��sWL��yX�\7���¹�1�y���� ��T/i|�s^�>	�"�)̠ɣW2A�3:��b*\��`@�Qn��{O�c)gWt^�Ez]	ޱDr@�H���o�Q2R5�6f����Q�d����(#�[��"ѝ/cR#�|�T�>��A���I�7t�(��n�8M��C$=t@�q��_�Z��j2,��9tԍŚ���#�������V�H�����J�
�j��g�z�@D��)Tl��h?��J�~�1H�ϝ��ye��i"gV#�&%���y�SO���U�� S��38jER'��9��U�^����v��y�n���g��cWb�f�ɚ4�}ٖf������g��n��2�v?�La�� -���N�/�Y��D�7f.e����g�㤁W�8�U�������V�x�7I�,���<I5�E�WL�1�ו�p��^�x�eF��f�Z/������
��P�ހo��Y:0�3!rS���u�{���� �z=z�N~I�m�G1�Z�$���\׺e &���L��A��������)U�w:2���B_^��t6���A��^��Х��ي��v[�,L!�߁C�Y�]xN9�p�Z��i�=���
�9$a�}�-�O��k�~
;�Nf)J]9^)�AZ{�5h֟ȃ��^Z�ؿ�ӓVz9��O7�m�o��Ο�ǐE�=#�ރ��ՠFݺ=%j�a��.�VRy;3e�΃���bF�-(o(�]%@�̓$&R���H����m6�*"�c����Y��l����>� 'X�J��DN;G=�$\ze��zNPW��R���J+�B\�X '�Y� �1�:����}���T�,1�#=3E�ퟑm0Պ)[�Z�u3HlB�C�� zż���u߃2�b.#�4��sa��N@2-��� r�%��.i}2L�:^�_^%�ͦ��k��%�u���	��Zq�i��7���~��t'@�6�!T��ނ��Ff�/6 ���c�i[���5
L��2��E��S��=&�����?�n��x�^��^��
��qpV�B�P�;ĉ�����"`��u�ݵ�cz���LN��~���o�WfE���`�����s�W����%�)������B>�F����r)�%�#P���ad��O7����~|��ز�-��LAQ��LS���si��<� ��m����ŗ�.���O۷oǃ<�#DBV��(��(���o����s��z5v_�\��Q"Fc�Z����[M��c7UJB�ȵ�7��Gp��c�]@/[Fi��r��<�R�8���@��ݒ����-8r�Q|��c�%����b)[l�����C���@%o�f��99)n��W��%Ge�������q�����xC�T���X��>7�����)�f��%�cd�UJ�LNM����t�j�dw*-�h���v��G�^���
�h4[�f\(�z�*,_6�n��L�y��xp�&f;H*^2���A���O�����o����|�aɌ?3Q
�S��tȈ�f�l*G<H��\��[LG0�����1��0���_o����`J��"�E,�9�ЮA~_�J<��B;�hw�`����9�e��}�R^��tzb~Ԯ���]���'1a�9�(P)�� �Vrd�����8<�4+�4_�{�C��j6R�����93�`�N�:r@��)8e�T]V��-[�8�ק �z5A��:�n�"h�_�P*���;N5ߠ(�P6Jփ'��nkri'��%9`�I{M�E�9����L���	����r���!�}1�R��qw���IK'�nFz�-)Pf A�V�<9��fL�X%)A�)ٴX�,�_�����,z䌏� '�d�;�e���&z6c����� &@��H�����V�ؓ{'��	�W�,1��tP��@'��!��y�Z���rt<�� ��&0%D�DNQ}'$3>��>�tXŲ
��7��<���{�����$F�T���]�s�ڦ��<~s�mXw�FLT;@~�,�$�+�#�-h�T@���;`��lqU����6�5���M� �kF��V�wWI��dE0J�@HU8�P�S��R1��K�2
д�1���T���]����@�)�D�%����gK*Q��S'�\ګc��R���,g�5'���_��2�c��ڵ�,�@S�ڈ�~K�?A�}H�t��䔮I|&��E1����{D�=SrU���8�F�=6J�/"��y�����Nt���̓_���w&��L����G��\qAp�_�n�g+~r�-xbK��0�~V���ˁ�Oc�^�|l�/Rb�/��Y�g�-q�	��Y��٪���:.n1R��G��m��o�(1�G�Y<��-��o/�kԹ�Z�0?�J�k�}�~$_BT���I8dJ�wl:I���9��T-���Xcm�
�є]IB��qb�
Ql�H�.�ǼR�*Y)m6a�b��䶐b@I��@i�J�J��ƢI(�v�K��+�b~�=�}��ےd`ڥ3�ɫe-�8s�͏�y�:]��cʶ�|�,�T*�6Uⰵ�H�JTn'��-4�>�֞bI*�)Μ�Q3��{�|R$�K�������6ИF����������;`�q{���j�@�#�UK���-�&��"��\�S�r�Mx�N�W/�+V��;b��4C7��)���r��]z3���!L��q%\��.�c�����|�W)L`���s��ׯ��/�g���B������h,L�T̢RɣR��Mg��3N}�e��F"�K, 	�e�|������eՔ�^}��cJ����6<�������_���bؚ�Eʛ���cӦ'�b�r��T.�A� gN�W5��bZF�D�x�	(���Gq�arb>�w�UG ���i�|��Gq��GQ���Ӂ�"�4��S���J��r��5��:p����s	+�~$FiT��п&�f���*�m*%F��� n��,�G?��P�[(��<����~��o!104$�4_ ��C�VEuf��Кĉ����O0���J�7ڸe�����06>�ݖ/����/`��mRQ����o�˰b�r���Wظ�i�d#����NuP��ޅ�}*E]����6���7��Gv`��G�4���a����lafb�'� �	���c�O^�ݗ��j��<���xq��e�i
��VШ7�`�Z�Dy�`k�r7���ˢT*a|lÕ"ȝH�3S����__r�zt:��˃HY�������Y�}4p�y`
0	L�<Ϫ[��x3)ǆ���#ckB�^(�L����N��v�*����c:0���,�l�^��MR�)ZU�Ut�u��Ҁ���{Ti[�������,� 0M	0���M�`ə�t��{Li��S���똓�ؚB&��^�3��J%aodȀɻ��̀�C��>vA�9v�k��DJ�x`�-�TF���&��W����H��cIL���	Ͱ��b����V:�LG�h�� =�%彴6+z�����tUr�|�j�7���[�H��`��o�$�tn����W8~v�mFj
�֪�?�d�;J��q5J�� �	<�@ڈ�c�Ws/q��$���&sѺ�V�J?��'&��n��X�V����C�2��=�$
9�����v>�\wG�;�u�)8����d�e���4�~M]4�n��)\��~l|���Z��H��iΏ��X.��e�`�E�H���:~�щc=`Q��n=z0	Le='����5�1����ji�9�����$+f
��GR��$�u����dr���uz���3�&䵱�P�@\ژ�Aj��kJi/#y��es|�t%.s������1Ťp=a~( *z!o�(i <.Ժ��[Ljg\�*a��J��+1��O&�N�n�DD���rM�u�K>����n�fu
��,
�&�:d/����pΩ�`���I< d�#�k|����l?��6�|��m���kd�!�;��=��Z�9�f���l|�*���o�J�VI!����M�0.�[�������{E��,�N�z�Z�VpYT07�2��亰^�H����[O�K��|_&�W�O�S�q���Jmr=ʙ'�ؘ0��Ehu#d�,p����M��	�w�E�~��糷8�v�^s�����1??���s���Nq���B�������9�-#R���kw��'c�hn��0�мHk��Xb`�Q�C��a�S�֛ij��J�3;Ȋ)�l�|i���:�(��]tLi8��L�"#�gu��Y[���+1�*��`�3�E�6ҭY�1��Eo`:�\kQ-��b�q[����*�x�}0��E��-oX#�� �����&�{�I���1#���*���i_��SNM{Vjm�[�]��_���-]� ��{�\~闱�J������)|�kW�����ȥC����ΣU������2��&�}���ğ} {�\�i.�<�o�m÷~p5��
:=������MY�|���ؼ�~tk;��|�|��g?�A�i����,Z���z�d�D�|��� jn���|����x|���ف���O�S���Fp@��~���q=�t�E+�+E����w�O��9� ���j����F�ſ��Z����W�c��.H�)'Ml�K�6�B���?q���`�q\������}��t�^����n��tR���[�y��I�ZsS;���8���/Z�m�ɦ�Ҩ�[���Q�7q��b�U+�ly~��f�v�b����a����df������?�;x���Jǳ}\�w��"F+y���>?�B���-�k�6�,t�/apt##C��_ڊ���C:���眀ϲb:���ϲtp�-������+
A�z�U�m�r�zs�p�V8fgg1?_Eu����y���vT�	e{�Qx�9gb钊=4'���v���6t�d�*R1�ҩ9�c0D�G���Ty�����-ظ�M��t�%cH�
��y����Y��)��6�
.�@�� �D9./�RXDa�I�x���,�vK*��f�&��%���RW_���>���saE��}G`�s`J)��fO�����Yܷ	]�R�F�EC卍V�D���fZ �����U	-L,�k�a���.���	���H�s����iF����j�X=p%����O�Q`B�v��e�t(��3宵l��}&bg�I�%o$Z3��(U�NU�Ǚ��K�P�����.Wk	��	M�4ٱ�L�L/U���%���&F&I�gLF�m����.���?��>c��Լ$	8��D��+(�q��E ��&�R�2�qF^)�Ka���n��@��tgc� o<q�u��8h�*bL!t��e���a���S/T�����=�<�'[QF��IE�Z�S�� �*��݋@׋W����㘋���;��A�!*!ܵ6I��W�U���P�`v����{z�>�IB:P��BP@�,��xA��E���J�w� � $�ғ�$�O?g�s�ϻ���ޓ��>��K�̜���߷����]��������M�0JbL��SqWvE���a`�/�!2~H
u�Se����sLT]1���4���3�&#�b�(eB�Cb��>�6,ڂN����V��,�H��t.��9M��1Qc	�J£=�+�R▎�����S�,4`��0`&`��\ӊ[N�� �w�3>{.���S�<H*"Y���%x�"����:2�2vݡ's(>r��������^qn���_�?���;��g�nK�x�(�S&�)Q&���X�+�l�x���W�^31Wl����x�@�e����U!iϳ�#[s�3�Z�^U�k���X�⃋s�%�{���_�q�ݡ��jXd�`ۣa`�_��wyr!'j���\Ե�{5���܁�p��tG�*��l�?/
;�]�`�K5d~D5�8̟�o~�hL�en�ܘǝO/�{�ET�T.�g1����+��')D��*u��<ػ*WO ��&�G�$�R��NŢh'0��Q�W�ȗ�	3��w�O��p[�D`*����Q�
0e>���t�2�bt)j+#@��\]��Sg�T/��h��:�y�}�p������6[UD�|c����1^(cz��O§] =�"��0�+��O=�$�=���9�==zm��������a���}�ݿ�[<Ԫ���CÜ��檋�Z<f���ˆq�����$�Y�j%�"Ut�(��ZF�QB[6�������?8̳`���9t�n{d=���!�"94[L���!�k�%r��\*��0��H��Y��<���W�IS\Y@AEQw��Y�\��/��B���O>����xw�*d��%��O~�C�bL�uಛ^��,�X5�J#�d&�\{FGd��T2�x��:Z���0��Wb��=�݅���9_�-,J�5N.���B�_�$^,$�_Z�W\sV�Y�}섋~v��+��%��o .��v��t �(��R���F&��g36:�᭛Q�oE��;x����0�+����\Q�9E9��b�u�˴C�D�fP�*~��Ru`��͸��W�{�G�8*ŌcO8���/0��M�)!שׂ��>%�th��D�]�]���@�VŖ�k04���>w�A8��/az�J�����˱a�f���b������A6�	F@89#��	��U�Ul�߆G�7z�I���/�퐏�_��G���te��1e��y^zk+��Hy�$ɤ$<,yH˼+ח&xG�r+5&ղJ��j��vJ�cr�!Xe� �ɞ��0��b�|^SJ�S���=p�I�=�&C�|��� $��؈_G�3mku�Si�:�1%0e�� ���ʼ*PR`o�� �J�%�i���������B�B��s�(vt�(��9���1h��V�/~r�g�c�����Ie�*mG�%2� �xQ�0ө7�
Lr� �J�ke5[�$+��s�BpJyQ��F�6����)�����`�P�����!��/�cA7�G�p��Ѩ�%
�ܙcI�������%Q2���4�\�
�.dTL"�1|`%�����P�%���ο Յ�b�Ģ�ϰۊ�bVb�U�]r茐��RS5IP)�0��Ǔ^o��j�6F�ێ�������v5ꓖ I��}��DS������o�����EԢY���1$SmR���[$�
 Tr6,2Y���ΈR�ϑ�H`�=�^���o�!䞟�.���:6�= 呄��a����pA59����1�*���O�m�m�eױ��d�_]��]¬��lՄ��{)hO�2�,�}��lN�����q5_T :1�Hˀc#C�4��5�5���r����8�
t������58Ӝ�q+?�|$d�=�o ޞ�z�: ��ة�y�v3s��[ m3u�i{�=���!$y��<��٣q�~;�3�?�iqS5��T��+op�?�3��A-օV"'Ψr�,��S��'��:��Pן�����a�ͧ�'�q���~y��&��@|.��\���KFu�3�΋��tSڏ4�����fCN��״�Z)(�R��3��Da���臻��τ�>�H'I��M�����ce�l���mv�iv�/�;�Î�*��q
��K΁�8���|����X���?��*^zg %$d�)�C ���Q�E�@�E�1�<wEʛH �ކh�*d��.O��!�0�PE����2M"�ՉdWV橒1U�	;Sc*f��){Lɘ���F�'�H���KKo2_W�5t��QY�~0����X|y�2.�eL�ӫn�=�"��yً̙3��YeL�
xVm����~�)��⒟~�}���5�k4t����t��U�����A�r��%�q�c�~�Ř9M��W��_݉Uk�8_ú    IDAT�d��hT�HԱ����sw�Eƛ��1�ς]�����K�3����o[K�7����^�8+_���A�f�c�-�a6`�ޛ�E�{�������k�؊�C���>g"0u�C+����U7��2�����q?.��jl݆�S:�_�?�7�����Y���2�ײ�6����ȶe��M����T�(�����=��$��?�N3�dQ�5�A���^��{>����;B�,5ƪ�u�>��n �J�� �w� Sm3 )@ֿm	�F`z�5��#hƺK$��d�N'�����FԊ�@u�<t���31�SM���s���9I��	�^p9�J<T��>ء�n��	���_`d`3"�����p�?���6��n 0}�-و�16�g�3��ݝ�W�شn%��W#��>}0�=�d� 0��
|D]$��q!�����s@HG��K������^X�j��������Ǯ;ȹ�uL =�~������Aԣ��m�0MhW��T�2>�,��4K�D�O��o{;����c�L,�n����z�"��Z&�9��Lٷ*��5{�7~l��D�U��cZd3~E��]Huu"����8"���#���+p��Byx\Ws/��`��4`*IF�d��綤A6���Z�ʏe_X�������렿?x�fq�k5����?�QQ���YǨ
pФ�U���&�KL�bq�9e�f�q�U3���^K���#8m���J�\
t9���<K*0Y�X�zq���36fv䳨�*v�[�b&g�_��@}�5�ǒZP� NEV�{E�N�f��S�B)�川���!r5���m�P��r�Q�B����>=J4Y���AQ�nG�%�_��R�4(+H���;��2n��W�/A5DCY�Z��V���h?2�"��{N��Q���ӤȬ2E�_�:��QCy���������n�P��F2�D��XRzH���4�)�z'�b2fL�>�`t��_.�L~$�����v}wz.����%H��vg����م�]S>AbEc{�]B͘�f5���Nt
���iL�~'�v�B���z�'hk��o
L�S�iťhh#�\���qE�c��Z�0dǤs�6u�$�����l��gw�^fb@�ۍ}���4�ɖs�ُS�8��[
Z�,��������@�c;�k�T�ݝ��!�c��2��s���
�Ԥ��H?�����.�|�8��C1�[��5>�����/BX����Eobk>�D��`��n��eć��aͷ�V��$~I#�#8 ꌵ4�)@�àSX�GZu�v�nb�S�n�k��S�/=��6���ĩ:��ǔ�����)��̫���]����=��]���hq۩�¢�[�+���s/�]�RA�c� E0*�Ҹ����"�;b?|����h��W��"��D%�`ڊ�:�-��=�¢HG�h������Q�Qd͓�`KW�S/�\�F-����lL�ã(���\,#M���[\y[�x0wލ	��Yg~)o�b^̏8�/�S�yp<s-+깂���eԕ�j��A�ZE|l"�atE�
L�cj�4(W�щD�2�+����{��/c:wf���I8�=9�U.�M���k�����y(.:�E���^8XJ���.�?�M�!��z��o|	7����Q,ԐJr�c��v�횋1c��Y�,^:��/��+ �kC��G[���?�/N<� �g��bG��\.�?�-@�`�G�/}�u���g�~��T��Mf���Ec�ؗՖ��8�	+_Q̏Ș���S�2��3W�2�hO�+���m8�J '��7"1�E�|.��F���c���w�>�}h��k;\~��E���e��2ꎘN"�Q���I�(���x��������]�p�%?ļ�9�v�IR�O'�q@��t�-���X���_u=/}[ۣ?�A����3I�L	�W���Q,Y>�f�S$�dRd��ZÃ�"���p�{��9�;���"7�����=�p�3�_���o &���^��=�'x��wO�p�_����4L��=T�+�#ӥ��F�Y�N�ƴ^�0�	o_<�#��Y'cf��@g2��İ�S���g��4�!�m�����7�|*�*>��}���]�O�� s,l~�˻�x�Vx���NaL�J�=�dV AP��AWeAz��U`JW�Z,�dO�Hy�'�b�/
�a���h��Q��GԹD#�uv�S$�g��5�AIG�z5�n��r��H<�LW7�=���+F�;�_��럀S�Kz-TG��� زD��qʃRܰ����3.j�$_� v�!ĬX���9�\Uu7m��]ф�����<���-qe�b�@�1�.���B�V&Ju~�dQ>+&�4��f��a�T��QV�;弌���S�_�r�j�r]$>�Ϣʂdq�%ZZ�?��9�	rh�2��j��k ��i=�N~f����\R..���_�$��qc�5�����$�f�#L��/���q���_(��*:Y���V$KE8���Dʀ��q0Y�$�	z&��G��+��>ޏ�XG}t/�����ˎmR|6ѱ����0���--<��b<��K�0�G+�!n���sI\vE~�4=+tϨ��DVhq�KĐ�Ʉ�m��)
�5|O���$W�Q��;NA��`�^�������/�%޺�p
tFЊ[&�u�$���%����I��`qU��:��aq.ڡ^=��^�Q%@�y݇sc�l5���
XT��!���#���Y�A�\y����c4Y���A��|/eU"���#�oVt�*l�\��a׳?��ӟИ�3t!U>e���2�Y��uͲ��!���2.�����d�O�a���c�ێ���9ڙ���6S�x詷p˽/`�`�h�XJ�'��!��3G
��+�i���&��'&FI�0a��롶;�]�v�gn'�p�6�@A��{��܋�����{ۺ�A�~��ql:㼸��S�D��O՚_��/m��V�D�?O�J�L�E��	�窓�k���e�;G���2��/��V�]�G�p�6k �(b�=��+'��v�ko�݊����� �A�
���:�f�՘� �l4�vƊJ��L0�]��vE)/͏�q�6����44���hK$�7PEid�b�xٮ.�U�ȉe$`��'E{��ժ���j5Q.���dM��C�0M�g�[qJr?�O�,>6dL0=���1uj��L�x�h5[��j���=?��B;N��wN�,�>t����4�K�x�������O��Md�S���puԗhȱ#�h��K����:p��Kpݍ�bÆ2����<��<��m�u�^�i�u�'��%���7�`�抰^����&>{�!8�+�<V⽉5}_�E&o|`C%����q��bö*Z�vD��K��*}Ԅ6��b�@[�=���|�sh����LOS`j���|r�!+�q����|�� �7�^��sl�-�3g���G��Ȇ"Q���W��[�0�`�9���?����"��i�����q�o��Ȣ�J �� ��P9�(���8L��faX̏�ک����?3���T�Z��?�g�Y������2�XC_,�@:�EwO��v!���S(�[*�g^ţO=�R�C.�1G}??�,t��2�_��+65�[ƴ�6j�� 2<D`�	��0��A���p�g��
2�)�:�2��V�'���d��UP��S�[mE��{������?%,�7O�2N?�����9�Q����?��4��۪�����Ӎήv�
yl�_�����`_9�0���0���T���+f���LTJ�W���$�,r������p�_oD�T�A������7��/�s_��\|'^}g^,�x:�TVg�Jo$:���.�=���+���0Z�k��G���q�M�#Z&���8G9��qaL��r4/b����ڐ�G�1�h�}y�&3���c��)M�!�مܤI�٫��j
�����b�So���/")�QT� �\P]���xش$����lH���2��1 �h1@[��3��3���s���&x�K���eبb,�4M
��ea3%94)���GE��{^bz�D����'�L�d�q�D�dI�:��W먖k(��U\��v+0�B���������ɢ,Q�= ?oف�:/�=�vd�"�&,A�)��*��b�CRK�Y�ҽ4��I�\8�1�gy�\�Y�0ĀJ+��A�P��]p����۵L8#}X����ЩCp��k)ۧ�R�9�"����LVΟ�jo�z]��<����K��}�/�S��T��E 1�����]�_����(���	E/	��M�Mf�r�?2�v�3m���k�ͭ��&�Y��
���9)�((ܘ����Q��xiA���� �z�����O���@�ܓ@��RJ}>��:`���\s����G�<2��歿/�$��	 T��.�¼�g��T�6�=�a`�k��˙ꇖ��~D1�ј����|�sP�(�q4/����kg.�I}NU���{����z���T�O�Ǚ��);l{Rڟ\QØ�	���\B��:���g�e�(@q��?�i�"150;���}��/G�顒Fqd �c޴N��q8�����U��u*+�k+&yi���f�_s'��܂F��eЌ&��sX��A[��S$����l���
=��uj#��ý��}�_ۀ��f!�¹��=s_�Cv�Ӻ����1׮�E���SW�җQՉ=)I�Bh�c�)�CZ鬀a8e��Z��kg�v�^f�u�erD[&g��1��<����h��<;e�WA:�a��̘ڇ�-CX70��z�d�tF�ڵ(���N	*W��F�X9��j�1s�5D���:1ƴ��i��\K �9�VzLI$j*#� kJ)o,��)qӤ�1�`{��>������kj����h��jo��y���|K�|��OTz��o5���`u��Y��θ*I�pZcS�������|��ʜ}��7>��>��/�%0����٧��i'�~�%C�P.�3=`ݻZ񉇕K �Y�e�G3��^���/.^�f3-���t��,n��bL�ѷ�ƥ���һ�vsY��6��� >�����/��ݜce��^�P��Ӻi�ܒ�����z���8�dK�%�^��؇8���y[�ě"�xwًh�p��Oą?;m"W��I��� ��\
�qnۊ=x?֭~�j�Bm���i�]���ǁ�0�{'#��a��2���O���$!�?{2~{�Oq�{�#C���]�0�xa�ӄ$��2�1�B\*$<(�?VB�4���F,ة�^�]�8=-�V9;��7���_�6J�4�M#�� �"�QA�8�Fc(U<l.`p��M���Y�T����cť�'��d��ž�7��p��b�;��$�ŠGV�n����Qo�G�0�Xm�$0��L��,��L[��M�6c||]�b��Fn�6tuvv���)s:��+.���-�tǃ����P,�_����g1��3k��".��[��ҕ#o!�փ��nI�8�;?�k��;]��?{N>�`t���FX��}a+��$/�,��)�c�*�(��-�|�����c|��}����N��*᳂ͦ<p΅w�����(0e�V�eW(�d�W�]bN����T<O�7��p�ʫ�[��28Z�i�V���*�2��4ڻ���>`Li�d������qmJ��Q��4�c�����G�,�� T���p4`��Ș��Y("NI���U
º�r^68�VN���R�p�:e��@vWMw���±�?��u�R�V�5�$) rzp۵J�_�����$�VM��K�M��P&��dJ��`�)�ܲ�x�<_��o�Sv��*8�ٴ5:R��5�/�P�{��tʎ=�%둘��2��PX�Iդ`c��9 |��K&�"��W�Y����l n�����DL��1IN������g�\�?	���mC�~��ib>+�������l��i	�d)Aq�q���

�[�j�c�]&�K�����v�ZC܈���j:��xz�J\��XݟG�K �lC,�C,��0���R���v�hK匑
7d%�8ဟ��K��+x�u�������j}�W
�^+���,m��{�*�t��Oa��:\�� f����|�FCfWJ�b�.��|�4��F�(�)��K�9)R嵱�"%�s�$����WK&�92E�$�n��@A�������ZP�Ťh�dR�.��P���6#4<?� � )�>���e�]{�\K��I!M�T^͏@M�ieX�ೆ�U�.^c���N��M�d5����I�X�v��+(v�����Hߨ�ѨQ-�+lCg��}�|��O`���B���>I��4�{�����4��<*{��NԣY9�x~���Wr�2�Y>��:̞��:ޝ��������K�B���#��]�2{���l@3�ط�gXؕ��'��6"5ƒ܈`NUI�7�Y�-�EŠ��z���)���(�%��A��}���&�&_�{N������d�n����m���9�\�v���mq1N��Ge�k���dV���mH_��%D��%+2�2<��cJ�t� �	~�!)�0�f��e��ǔ�)�����4}�0e�i�3'�� S�Ċ�6��9�TJ��J�)�5k�S���m�r�N��L����,t	O,��*f�:�����/s��zAM�(r����
�U7?���$��%̞ރ3O;	9�4�U�5����n)�i'���e�|s'7�^:H3����u	�t��]g�wݷ���6m�K"P��ym��0��p��-݆s֑1���yU�a����׾�3&'D�,f8~�)m [��X�|�y�M��|�Z�e�I�t���^@�`�E�X���L��6���_D�8(�b.��>0�"�c�=�%/��g�Ba�3W���Ȥ�2k���T�bpxc�<v�cv�u/����X�5����wX��{�s������?�G��E����~~�}x��5�62�#)4<�n��	�)�U��@�VD�4���z�>�����;#+�V���z�-\w���{�}��; �K�}�꧀V�U&�*"(WX�a�_�&��6�}o��8��(~� ���1���.��n������h�Ǘ'S��5P*�0>��R�� �:t7���3Н��hK*<O<�$���D���ϣR(He*��a�]v����}�&i��9����\v�����|x{��t�mx�����'>�s�<��j�SC�7��۞�k�-����� ���#tad+6�z��:�~�8��}Е$05�[?��R)�u����/�[�'��&"$՗��^�+��w��FG�q�G�`�ô��}@�S�݉%˷�C3G�$3i)T86����4B`��H�Ԑ�ɮĽ���Ϫ�@���=h0~Oվ���<���	�\
E�(�e�����@{η'����1QN'H�ڨ�B�BQ��d	l'��)Zd���@�,����H�B^��V[I�t��iq�GQi.����H��jk�[��.c<x|�P�]i�VIZP8�K��z�a�+��:�}0 j��}��Y2!��֫.�^����v�������|\��ac��A&��T$9o-�g��1�5[��0)�N&��}O���G�������
��l�4�P)���APܱf��93*΢����v���)�C�@���Y��W9�g��ٚ9	��R��p�*�*�c	�ȥ�=X
�ڳ)�,��[o��hlTKh���� �w>�����{NF��4�Kt�-`��n��	<��[m���HI;K2�U ls�E�n�0�J�ʴ/>S��Swϔ	�1_{6�i��
�0��'Ųl���b������gt�	 �}�yHZ���@�HBWi�W�������W�W��Ep�5P)�իH9��?�ro�,ȹ�"ߓ�]*���_���ceB���꒫y���<'ƲT�*��Ȯ��$���q&��	"�eQNSF����.�ٌ�|}���l��|������K��F�g�/�8hy�s���b�1	���9��8
�,�t1Ɗv��v�!�s}�Z�V�    IDAT��\��٬��E��Z~r�*z�|��ɏ��wV3G9�l_�Q󲨐k��;��
�{r��q�"q�Z�S�/"�1�msT����H�q�b��9b�}�P�ˏg�o��7�74ܺ}��_�a`(g��'���{�`/Z[�/�WGh9��,��W��3+�ʞg�%e�"[Vy5�d��ITnMb�<�aߔ�p\�RX���ד�!�`X��Xq�YL�#�Fk�R`JbK��/��
�B���*+��!.R�����3�J#���GI��uZ�P`��s�Q����6^�8R'i`�4�݆O'w�Iև��&�H�먎�I1�R^o��ڳ����Zx�@ aE)/��5N|(�l��4�mCL�&-�:�f�cj��y�2��DƔ�X(��5��~�����НP���ʘ�_��/���	\ǣ/aΌ^������CvG&�����G���o�������-����������<�P�����~��U?]�r��P��,+|��Z]Í�.½,��h�H��v���_��&�eUj��\��;�a�&/�r�h]�I�4w*�1
4Q*kOD����Z������a4߀�{Rm��q(.�+Q#΍T&G*D�P�DW{
����β����k_8�<���2-�>���V㟷݁�a��HL�܃��s�-7��{�z�Bk׭��o���#%����r�(�X�26oA4��;��e����w�A$��_�G����.<��zԚ�*O�*�hq�q{31Ɣ5�Z^i���yV���ˬ��Bj��f�<��8���1e����s���^�3�7�+M���t�[��tVȚ#����L���.�9
J�_xk���X��"}Lb*i!�c�f�T��14Ky��[��#���?=U��µJ�2n��mX��3�7w6�^�X�D���1c&�(k�'P��0::����r�A`���I�Ձ[�W_w>���q�����LCL���MU�������q���ȶw�or/�R��<>�m�C_��IG�|OtS	�,(�eI���+��;�����T�%0r������^�| ;̙�H"-}��ʸ���#�/��}� �S1kZ�LY�a���܆%+��� �mG�-`L+�)Ѥ7�v��)�&?���G`j�Ҫ�r��n���@5_D�Nq���/`�ɞe]�!�J"�J�s���H�&�i�P@�P�ĉ�4�q5��1-d�(IfN�������sL�����U( )=�����s(��Q�,�Vt�@�O�����S�O�����i�$'�5i�J�h)����a2����^��&z���א�P�d��!_[�)|��������(FS$��D�9��*0�5��gʂH�����.��������ɵg�\X}|i�
K�����7u,�~.�?*�C��!�S�Qe�$10�HϞ�Qb���o�R���!ÀX�γ����&K�%�V��r���W�G��$'��Ϻ}���>��������^X��$k�������,vUH�]G*��*JÛ�i��ȃv�7�|��L#+�`�~8��_g�\��m��+��K���h��HdH��'2*iff Ed�f��ٱ��A�@ ��n�\��۱�Bj����E���}�0#��Aem.YT9k��=r��a�A��P���	�雞���Z@%�V�P��F��z�,N��Z��jy�O��gj�d�Xg{�l}����jC_o�(�R���Mq��������6H�gU,ʥ����DZ�y\�tp���(�GGQ圹���F�J.�Tf��>S)��U��<�A,��eٶ�J4�H˸ο�`w���*����4{f�Lu��^h�M�|�������-N��*�󾱙]a�ˇ��w�x���-&!A����`�r�L�B��ɒ@��A�$�r������Ge���'�ۡ%!�)T�n�C��g��[��u�5 ��Ţs�$A��A� 曃��t��u���� f��u�\ ��#�f�_Y�P�c����/+"(���q*7&Z%l��B��ܘ�6eD�
c��x�=�ČQi�h��Z bN q&�9�����t�Y4A`�muF���KdIT4h�F�S4��b�',.4����ĀP�+V`t�]۞���J���m�l�Z9䨬_��P:%>/M
�d�0��2��o�φR�q���|>�z<�G����K��)n�f�&��0�Qt$U�[G����
K"Cƴ=�F"*ƕ�
����'()/��
E�l;��\0ukZ�B]�6�U��V�:�'�Gq�
ېk������?��bc��9)�)��x������h��u㌯����ل�ԭ����>�8�9�`\p�Y���\�N�Ĺ���vrw��\L+Dlv��HI6��5���p�/��1ov����&�x��~\��۰qK]fJ��u�������/��^�,�M	���t�3�\�x�L;:��H���7IB=�p��ڒn�3����)}(oº��#�2N<���{_��pbF�lb��{�qL���'>v���q,T��E� pc7�3?��x詗��X�v@��ө�{>.��Y�k�IHҙ��Aέ�'^Y��F�h
�lN��	(���1�b�LQ��Z~3v߱�:�;�?#�(>;�a#�Ν�{�$v����GQ��_�ePm4�X�z�|�]x�����#B�O~l��S���s���|�����۱q�$h��u�;�-�Z,�26�Dc�:bO\p�Wѕ�D[�$0iX�tFG����T*���!���=",,���NE҈&�oDp�#��?�9p_���o�7AƔI\oo��Ϸ-�L#h��Cߤ>I4,��Q�(mű�-�WO<S���\L�mۊr!���RI�?����VC�^G���]=H�1\�t�\q�mxk�{�pȇ?���U̚��)�2����ߊ�+�!�t[��%+울>��(8��-�a*��-V͙�6[2.&���T�<��i����=G��յV(��*^�,���.$ڳ@�9���}��3�X��XB�r�RY�,�L�'���J�����b��e��6�8T�!��V�(�G�~@'�PϊH���T�Ԥ�
<c���X�ă�﫰d\v�|�R/l�2������&��3#c�E�mɸ�;���g�&)TC$�^�����S��Q`+�C֓˸G=�E�gV'%��CΩ��Ei�C,O��U,&�r��r��
g�IB���s|4���{�E��g?����'�T�q��`�����ք�[&Uf;�҆;ai�{����G�@J�� �..��~N��y��_\���\~�c.�z$ZO�/532��x�ʴ��xAf�kЬ���G��cǩ9�����O��]br�g��P�>�M�ux~�\�#X���Z��V�d��2�d�d�C,���L}z+mL�.EKlm��B���  �C	`��O�]���'����{���~���ٸ-vL"��3���q��x�"�z���j� ���J!OM;�S	��&g7�HD�M%��$�ёÔI���8��DOw�{�eUI"����K?�����S��X����7]�wU!��b~Y������W�����7Wbd8�"ّ�'�t�����-�<��Ld���mkG���x�c7U=�'�X�I�I��ߐLr]�$��3i5��4�C3W5V:gX�3��{�� ̭Rk��IP$nɮHb�q��ZK���`��1{tem5P��Hy��0�kN?�3��9�ʹ����XZ��ԇǞߊ+o��Z3$~�t����)��~h�Za�ϧC@�m%']��vqϏw.-���OxS>ٞ�8�0���1�Z��Y�+���P�T�=�V^�rw���ŒF6�U��7-��b�\�ls㯜�.7*�a�5�,�?���W�ǖ�a8�3��!�<��Q�x	��Z�k���G_��r��A�R���d�,p���="#���@[zƥ݉9!D���W����ɘ�D�� ���@��S5���z6��4��Iۍ�pi|O"�юXG�x�gLyJ"�9��=�;FR�[/:Ɣ�K2�i���$�A�7��ʏ�Aɭ-�b��0N����_��w/�S[j�"�V��*N�����˯��#̞օӿ�,����&���<���D`�v�5_��	�3{2�R��Y2,���1q{d�/~�]�&c���S��!���M�EGA�^ҧ�ي�n�Gf6V+#�y�\��ڣE�RX��\|�mش��T�C*������V/�R Ɗ2�x؊���H�� ��@�)h��^U1�d�!f:j,a�au��SŌ�=���n�H���>�u2Q��h�z-,Z��&O�n��,����Ǝi`T�Y%yM��M,^��=�"�xq9�-_�d��d�3����cV�HH�P�li���K�D����x�H��̼��;�c��K���o�;��yӒ����*VM������%�\'oɎIݜ�C�t�#X�n��x����읂jyL@��sL�;��r+��_܄�_}'����I +�	r5:��VV`Z�#+⨃w��?<��15�F>�M7���0k�����O)5�5s�eh?���	������ށ�y�;����S��U"��?��4�\3��J��^����w|l��mزa�����]q�������gҪ��֮��ǌ�(9-,ר���i5��*�g��WV��WV�P�!�����Źg;L�ZOE ������w�|`*R^��ղ�Ti~d�b&u��	P�j`��1m�!U�6��3�
��C4�tR^a�(1`�SV��{�oK#�>o#L���~N�zLk����U�ɘ&'��U7�U@�נ�<���l)�e�i)[�:`]׷��Sc�$_"/P&T��^)tA ���n=3&�s G�А{'�s.��w��L�I�(L
��AYQ�4��K�'e�$&Y�ZF����n����i&�#�@�gN/���O�_��+��ZD}"�"˓���zCl�˕�z��M���R3�� ���!ЃA�]�
'X�,L�Ԁ)]���صDU?�#p��yM��]Z�/S0uN�~"�f�:eW�ky�3ӱϤ� ��m��>V �dN2cC��,���9�G @��ZΣQC�<�=���/�#�'n���(��⤸5�H�U���x�{	��5PAV�ܣ	�&�� ��	�&�
>TA�=��@�<5�pK�b����G0���_e��B��T�(ǹ����&�nM��ͤ&]Z�R`�ɻHR�[\�h2�b�(%�e�/�+���&C&CWG�����Ĥ�N̘1	ӧ�bR_z��1eRfN"3Su��@�l�ގ�a��]���![�~ﭲcvl8|m�[7��j,2�{lX�n�n��x^ڇ�^�C��6T�{����M-K{�UĘH�j���x:+�L[;��mR d�$��L��c�J���K]�5�	z�sZ/`�� �P��U٣1��	cB�bnU?W�s��}�jMVX���h9��^o�&�ʺ�ZMT��h��h���`��N|��#p�������aE$�w�w�u�٥�����ҲM��:�E(g�إ�WJ����9��-�^�GGG[B!����`V��r��	gB&oa`�Ԑ��x.���a�`A>b6��5A�'J6t��:j�qx�����?~f������[&��Ո�E���C2��O��4�H�,"�G�{?�.�Ⱥ�K�!�!K@+D�ԃ��lX!!$C7�mee#�\��B\=U�O̥ö�4"R@7\���X�o�Dƛf��X�|�|Ir2��]�u�K�Ep���,/�o�4NW^eL���2^��4ڞA+��:�T�L��D,"땭?����9$3rYQ��jB�I����͇����fM�^�Hih0uRމ;��-��Hx ���k�õ�apd;L�ķɘ~dWd��ŪuC��W��B���)S�ٙ�>�t2�W3��#un�s\$�bH=��)"r�HѴ����v����wĤ���B�hf��!<��"l��W�n;��ګ.��>��l.��������*R�vT�u4�MԼ���4�k�+'D-5��6j�f2��	��v�wMA���]�����Q�Eճ��fڔT�#ذf9"�q|��p�w>�����`T���'�Ğ��ys����1�Aj��a�,~�]���Kx��Ux}�DYt�g�ߞ����DjGg����e�a��!�	ԛ1drYu�ee��#�jp�T�伮F��f�s7.���;5ꏋ���h�T,K���!�&�K\��j&��֏�wWބ����nx��|���׎��y�`��Ӈ_�ﯺ�Ze����t*���b^%�DsG}x��_D�s��\k׮G�\���s����[gz�;�>�5i�Z<�PiŰ�wp韯�;+W�'���i�v&Soo(�O7=��W�`��L&+��]�cp`-�� >��4��'�������)�C�_=��c�s�=1o��&cR��$&)�z�@�E<��������52K+��
0=�{_��&g����ۛ����ߊe�Fь�ȴ!�ͪ	o�Ր�����]�\�HK؛�"!�)�̷U���ӛ��*0��(�!�\�Ӷ�N$(��(�Ԇ[K��h��`Z�T�K	"��t#=��TRf��1�1�X�S9��ʞ�ZP("�
���j2!���yJ���_d����P�
{Z|D:'�]�&Z�SZ��:���N������;	��٘�����Ā��%Xr2h�Z�x�8)�v�kQG�3ȜXO��qe�X���Ń'K�����L��"c�֔Q14E ��i�(�`�����$��-�EU�.� J$���g	�o>�E'�t,�|^��n�v9`��T4�4K~�>�/W(p�A��Ӏ�c<v���u�(
��s�2���s
օe���ԩ����[�D'�b��T]Q�@�=q��e�k�C�<���D+��k�$|��������EKJݵ�QR<7����;���o�G�K�X��c@M˳tβ��bVm�U��H�_¼�(Cw:�G,wL�猟 �dZͽ¿�5$e��0(U� ���d|���5���7�{&E4�*�����rɌnʨ�@�$R�(���0���6ӧ�a���c����6���9��'�v�{x٪I�ר%���{`�"$/�ul�ʀY@��t��P?�(��������k<P�@\o�𗄍����r�q���7�����UX�v36n����0�e�c�L��,�B"G�چT�]�h"�l{��$2�+p����AL��lM�s��'q�s_�7I��/On��y��V����gC���OA��Rw�캯]P�2�����Q��<�rW�Z	����!L�㘏�o~�8̞���f�[��D�8���w=��]�j��9�5�\`�u�eA�����.t��7���@����s��	[������/+0:`j���W�g���
����F�^�"E
�	�RD�2���$�7��'�����
OQ�~ϣh�ǰm��\�Dmh497�J��d0�V��R.�Yˣ+����ݘ>�[b���8֬ߊ�|�l/Z���O�[�����Z*���ݹ�L�+�8�y�7գ�\s$q�F�)����A<�7*���6A<]�|;�-���PT`*�2!��!2\5l�3��w����%�/�)0�W�R`L��!�A)�1�6�GZ���T\e�	���C(�fޟ� �f�G��[T�5S�H!_����78{�<�\sg�r�z����<���������<fO���_9�Jy[1��0��W���h��G�գ.�I��DBθDkS�t�J�C-���7'C<����d6�d��*�z5�1�x��F��e^n��R��O]v+M��6���܎[�2�"_*J2�N��-��̚އd"�u��X�f�n�3&a���b�=v�Z7m������Q�q�	5j�����ju��Yݝ9Ԫl\�."���O໧%R�H҇�j�x���q�g���g�mC�Ez6���c/7Zx��U��3�bɊ��v#�����3��q2�o�t0����O.�+7Qk%QkD�L�EFB'�.��[�&��rU��ܙi\��oc�YI�5֩a^K�y׮^m�T(�]�    IDAT�A���E)F�6�uv�\.�-���i3�g���~�|�cxv�҄���p�G�����y3�R�Q�	<��F\���P�e�Lw��q�aVG����Zy�� >y����/��\X(<xc�زe���ȤR&��:��I9��*���{��U���F����x������}p�O��s�%�{km���x��m(�(yk��H��V�0�u#b�(v�݁����͐���eo`ѳ�b�£0g�-�gO�"�5�J^�,߄�\{/]�r�6�� '@ؿ�|���S���Y�L�}'�X3�r3���P�l����6�gL2�,F�D��sLٓJ�ug"�w�&����ʥ�qcG8��P`Z�iY4<#�p3؉�Nu����Rb�T<�݅��^����UD�t@�ӝ���b�&*#㈖�H1��^X�.&)c��!j���(B~_J&�Ta[�SFH��-v1QR��b��Ș���8j�A�Fh���4Y�&_jޣ�QGJ��F�'��VC^\rEɓ�ЍL���:7M+�4��WOE�<��Q޿&��׫T%~�mL
/3�J!��K7�|�6P,UP��UҤ��<���.M�D����y��D3w���q���w=v�[:9���ڡ��
�1)���� p�i@])�+�怡r�)��������"���1��l����(�#�^�a���L;���a4ZkT��yyt���Ⱦ���/.�.�3�*�-0ڒ���5,Z�	���4Vm(�B?�KJEL�Q(Mo����S��& yn��CV!C��!��zb�W��Z_�w��튞�������/�󹹙vI�4���jJ����$��:�^Q���*"���<�8:rIL�ԅysf`���1w�LL��DwG
���N1�DH���Uk%���([#�2ë�i����&hi��T�u��q�����i���B&�B����/��Ek]b$W� ���1(�(�j�c�,_�o�܀��#�ad�ä V2]t^'��ʦ�a>G����s���\YG���&0��f��>W�u���7�9%I��Ѕ�
H~�C㝂��Ut��5�Xen���ؑ����#^	�H�ýx,>��T���m@��61E�v�;���Ex��i���}$�g�Øa�P�M�sB�~^�'��֓+�Xl��qQ�mL+BI���_D����r�R����ޕ�U.w43,1	�4Q)�Uˢ���j�qj�Yx�g7tu$�J[��ޞ��h����m��O���Vb�����ST�r-���T)�V�cF_
�?�@Q���+ �x��u�����ܫ���LYێ3F�Z�>V=��w�Ʒ�8_/����7RWr�#3a�X��O�1>G��G_�;�1�)���3&��QdI����4[�b1$�;�j�4�1�V�sS��(���ő�+�Q+���5�ކh{�DTS���D�0�M$�!@��rY��R�LƔR^z�����cJ��6Ds7YQ�:�� Ӭӯ�~t�*���Hy�J�����%��o�ah4�YS��S>�O��qZ�Ǳv�.���L+y	��R��jl�(�}V��`�����N�6W�
Ò�1��̐�N��	D*�mŸ�K�k�i����aZ������p���c��
R���������ߏ��1̝�����2n���X�n5~p���o����T��-��owb��[�������N�+���yW\�).�a����}ѕ�"?�o��[7�C.���v��P�t�ZR�dV���d�j���j<�l-�^����IGv ?poL��D,��;k��7?��c4�i���}
�Y@��ȉ���e6X����uGљ���#�~���̩4�IT�B�������GG-���ڲ9���I2�eho��ӧM�	'����v��U��K��+K�P���Ì.|��_�왓���q�P�籗q���c�A&�%r	<�P>�a�\@^^q�=�>�s��K�Nݫahp/��"֬~3gL��,7���(�J�h�d�d��V��T18^���X�X�5���V�b�]��{g����O�D�ʒ�q�?�{�P����4��4�&V�:FG��0��''p��O���\?��"��~�cX�����Lu�3sݥƞڲ���"I������>���j��P-0gf�:�s��G��1N�-`���K���14��J�l�T���H��.t���C�5J�f��xV�6ī#�0VM�����m4}�z�&�Gt�K�e$P�@F�Xb�UZu�#�NФll\����0M��J�i=�S���>U&tլ���Li��~
e������p�3�JyuV$��!˱dԆ&�u�W�:p:��i�R��]�_E�/�j\�ťO�U5Q�~[M�����Ru��*��F�gJ%^�l���%Dܯ�y�$+jd#�ȼp���h!}c
L%M�y(ڨ&���"���5:�� OʁUd�i�*=kbO�����������~/�S��z��s&��# x&��ֲ tMn�d�n>�&��kk���$�Uo���f�;��n���̎|s=^%usL�V��-�M�r��`��W�9�&gC�%(	h5Q���U9�wfO���'�3{��x	�����D��C��u���sxh��.%�E:MuHaN�n"e<���h9�2�#!|v��z$�a�Ic��ۙ���	乡�r2�$T���ξ�][��]����}��*��f��g)�^���%��
��1L�܁�w���޿�.�lO��S���߁P��6���� ���b�>"I�J�?�vl|�}��PH�0^���xXلϩV6�`�{���*.��Z�
��UL��|1�V�#y`ݦ*�xs5^^��ڈM[F�p^oF�d�/�D<�A<�B��َ1\�a�����[�T1F�^T���k̝(�v}�V�w�,���Uu{܁2���VPD	�$�d̍���=�2vsY5�]��j���@���7�9S�8�p��Б�}iЏ�8��{�p��S���{��k��T'Q˃�� @5Q*�2+�ȶ0UE8�隱��~�/!3܇��@N�s S��VsС�&)u㘔h�M΂(s!�
=�G�l���q�w��=��է�����RmX�rpۃ��'^E=҉Z#�dR����(}�(�ri�V	���ď�u\Ў�am�i�v�#��ObkhD�B�MOm%x_t6��?���v�S�~d]1���K\i��	�i(Ă/�L��$:5��	�"(��V����L�F�:ۦ�Huw *=��Wƚ��H��B6��y�1�}��j�9���d5?���`��<=��%R^z�D��Z
�)h�d�T��bj� ̀�
X�,��2έz՟c����S�>�l*�4��*ut� �|������1D)�6�y�	Xx�dLc�40��n��<��<�uZL.B��^�����h�o�Kt�������+0O�`�ߥt7j��ZbI���?��m�`.>��ōU�'"��/�p�o)�����n�*�en~z��q��E:J �|3��oF"��y�|���`�C.�|���w�[�A���d���� 'L���}'N�Z	YRE�4�h��D��=Iٍ̝�|���a�$��rP�1�?��Ï�Pi�����k�ṥ��(VZ�Ԑ�m�$�ՖBOW�ۻ08Z���1D�9�"%�Y���Lr��Ȩ���HӤ����2&w&1���l�8�x���^�	{��1m�dq�m��Ж�	(~��W���O`��iXx�1�=g.���.�y�M��4�f,���cJ_fL��I��Ĝi�X���l��`�] �HS!U)~�&hZD�0x4*y��X��\dS@&M�<F����C�U���V��t�-�F�Z��$e��tV���"Hd;�3e:��=�g�00T�ʵ���am)|�����;!�Py�[+�c�+Qi$�#�&8�DP�H��J��m���}����W��ч�&k�Zja������8�Oz!�L�,G��3w�D�*�R��uTo��=�z����7�X*"�p̑��'��铴�L`�b=p�/o��be��ڨH�\I_^J�M
�@M�_j�*�|��{ 0�^%0��_RP0�Pd�^�񂌋�j��2��HPZ��엫kQ	P���fP��*J,���DrR/��$�(��	�O�:E��k[kJ�)
%�ɘ�k;GQ�i�'Q�5eT�}A�0��Jh{�ӆ�,��O�]5��KƧh�&{�9ߌ�BAeZ9D�Y�Ҫ�Gc������$�Ji��f�0��V���
Өt8�1lR�уVf �O�ɕ�ߩ{d<�BR�ܒuT��;���|����J�|�c���'�tG�A�NPyf2�(��$�a�X���	�K�C�>e�����ukF�@�vo�Ӱ�>S&	��KC��pRr����:���t;9�v}�a�*j�c��������@�󕥩�H��̩�REu���>�ObO�Ґ� ������K�X^[>���{/-[-�]$;嬨7��c���HE�ʈXmF�׭x�!����a��`zP%��q�~h i1��ve$u���e4���4��j�>dR,���G��qi^y\b���6�2&�}�.�c�9�e�LL������{�KV�Y��r>uR��9'�4�@V�aP�4cb���w����u�w����
**�2� 2M*H�3��9��ʵw�����vU����yn���>�j�o߻޵޵r��~^�6�����m
���N(��ݫ���oۄ���iQw����0��Εڨe+��jOi\��{���G��X�P����Ѡ�^�̠jˣ���?�r�-U�CG�غc?^xi;����~�(�� H���I��$�Qq�餀�1^���R8'�m#i�Ƽ�����ć�#J��
L�=��+o�g�	�l���WF{�K��E�J2��4��aN�V3�q|䪋�痞��>��K���0�exa�8n���������A3��d�L^�}�Fpo�4ː�nj'�:�a߻�8�6@��a}'z�O���j�c�^6�)��Y�C`��v���SCu��p���+q�)3d�@Ƒ��0�����t]X�4ی�k�_l��x�	�>q�-��KS�A��f	�3��K��ϾW���U��"��{r���}�`�E�3H���ܲc.���k�$k���E3��7=�r>���vF`J?UQ���y���#�NK��L/��pY�w��1�O��VR/�ø�fq��1`Z�#�J��7�W^��Ű)$���iD���V�k�i$�Rgai`cq�����:C"~������1�4'������~~?&&+�1��g?q5.~��Z�5�6��?�#G&���H�i�7��Hͤm:)fA�D��S@3�E���	�%o,�}~?)�"rqY������ԡ,�-Vi��1�����C5x�Y��'<\x�|�KWcJ�u^$�g6����>��N=	�8o�f�J�׻���_a�*�R�)�,0�]d)�d�Y�-hi��
�~���.���i���0sz�9���X�|��_��t:�(&���${�5�h��:�-c��Zwe�Q��F�M�DO��e��h�g(�M�9S���{����]�#��6ЪO�Y�D"�F��YS&�#��N�y�l��f��K��l�x�/�֟��l�<}��غk�߼��N�ԇ�B�t�F]��̉�� b�3f�LiLn����N�d-q3Zr}�e�yqA~�	t8�D6���@�gc��A1����G�&qh��F�D'��ЌY�6g!�M4�e��� A)p4�t"�\"���*^$�t���|R�(�'����I3l\�o=�$R=�{�oF�<����q�{.�O,�8��Q\�ri�)��v/�~|y/������aN��Y��q�;��)kW �W����[qǽD"?�6%��^SR�Xen�t�e�V�%=s6܌YXqS$K�(*c* ��xL�OlZ�}�UwB`���)�4(����3nx"�2b!���H	�35�5:ks6	H��#1eA��O-c� ��AG̏�TƘ�j�i�� t�
�a�.,0��WPdyx�,�/��6�A��h{pQ�{�)Ff"���ۚ��lS��X�|	�Λ�ͦ�b���m�u2&��D
<��a˰�x)v�Zh�2Q������P�m��TN$�,��ф>p_�R	���r5��%��&�ަ�K;��4t�9i�"�4[ ;mK�f	f,�4ٍRT�؛�p2��<l�I�l�7�l��.��Q�����d7��@N$�&����Y��ũ�C��v��av�dx�%��G
.L��T��Y�=���#��*�V�O�̞�I�gJ�;�%����k.�[N�#&G"�6�_�58����/�mw?��vCty�6I��.L��\���̪Ƞ��{�i��
�uޞy>sV)�3�*�V~mfj�U��R�^I��ݣ��[6��j�|�%EB�k�^C�|\θ\���������u+�b�\L��@&�yM����]E��ױ?�������,۸&9ȱ��MJc�5��[�KTY���z���E=�_3U��|Xc4�_S�@��J����2�l��>���1m�Λ��3���b�Lͬ�؂]���¶�VLO�H�M3͎IR
i`|��J�ؼy�y�e���6/7�p�K�I���f���D��&#�d�eo#�>A�j�;�D8nb�v�@��l���w����њYF�Z��=�GV�
��x֮�>��l�<W}]T��ހ_�%�|���s��+߆�E �wFa�N�m������̋o���%<����)̩��5ܞ�V�mi�Y�W���i�I�gFB�E��F?�'K�����{�݂e�3&U:\��N}���G��6��n�Lt�<��K�c�~��D6
6�#����]M|���{����"�F���8h��k� ��+�n��l I�'�fF5���M��?�c�|�MǑ 	��Q�Ȉ�}�o��ʄ׆�rmmc�4�, ���Ɍi'N`j`��(f 0��i���<�)�8�e�J�BNrH��ak0��#�ϣ�\*i��F����K|���%�I�=k�)�)�^�-F�E�bm�z�R^Ψ�̡�o.S5p��%ɲ�M×�#��v܄Ǻ�1�$��3���R�0.& ~��O�Ƿ?��R������9.9���a&0W���ֈS�*����s&\���Z��_B���� ��Y����E)����C�}f~�E1]y�#�鯰�@M.V�)c`(�����q�e�EB��Qi7��Ň�{)�O�J�_��h�m��Љ�����Wp�o�A,1 ����Q��b,���K�@
=�"�F�[���	L��8���X0\~�j���ͪ���N��V#��@��������W�w��1'��%W��9ږJ�ʿ�R�_\�KJ�H��I�Koc7$E���q�Y�}̔r��ii�8ȦH���z,�я���J��~%R�Xy��@x E�Ǘ����B�ég��v,�-;�`��q+5�i��*�1a�cMJו%O�x4�n���jgZ b����{b��a�Q��n�Ѡ��Sr8y�L.��Kbp��ysg�����N�W�>�MϾ�F'�D�#3�p�cUqQ�yڲ�����'�{^���2�t�P�A��)W��X�E!E1���}2���8�=ǚ�3����.1��������G�H�F]���16���o�x-���{��
"��&W���B�\^'��ӆ�b�>P�aA h/�Z��6E�)�d�2�5�AJ/�,�QSeL�'��,q�T^"c�d��6��i&�� s����:�5j�%�q���6�6��y7lJyyf���HMB;�Žl5p/��S�{(!%�r�h�� 0MQ�k�y��V6(eL%{ј����|o,
[�J��@2xG�HG}������8�_�P����@+�.f������������h�dJ4t촪�2��ԁ4d�*��N�jLY��~�#e�m��_����:l Q�.�P���w�gb8�7"�Ùd�����8�43A[��X<��|�qx    IDAT4Z ��svL�0���>�Zq�%���Z�K��I!��"*�Ab��M7l1$���N 5N��g����i9iP��f['�n���D�:׮�^�S�)�r��LgZ��l�)T��gN6@���pb��~��rOL��=H��}�8|Ӫ��8���]����,�	qtd�βg�L`�
�y�K����pd�Gͣա1GI�!r��l1�]�K��U9��%{v讪�B���0|o!-m% �Y�^�d�ҨPĶW��0RVv�y��3g0erTT��j�Ĩ�)!�n ��1wZ?NY�ׯ���s1kZ3'*�OO���ck[�X���!
 �L��$0sP�4��y�q���0Y*����0Q�H����Ɲ[�R�?m+H3F*�����g#��������bhт9X�l/���"���˦�_�!�I"��!�� ���[_�Q|�I�%�)���Q@SE�����^�'�زc�yn�ev�;�������$�A
Q�3��C<%8�e�;�%����T[7*F��ffz��=q��N��K&�yvձԀ2kH'rvJ	����ݧ�f�Y�TM殗��:�`�*|��K�raV��I?ВR�����u���~�$��YT�:�~�Ɇ%S��7t��vnَ�gɎv�kh��:!�(s}��R`(�g�Ț��gD�Z�6�*��TX8d1�-��/�a�P���8g�4�hD�=xiȈQ�� p�u'�9j"�9��=�|	�t����	�"?4.UY�*ʓG�	&�a���K���eE~�9T�V}�7�ŷ|���N��r��L��+�*��6��8xK�cg��B���n�*��,���Ɍ��D�3����e�i���UWƔgl�d ��=�TS��!`
���r���:nK͏j��ۦB��2��T�n{�=.%b^���Om:��+���Q�� �c�9���f��!H����=��D٘p������/�/[�ń�=㹮l\L����Gq�/7�T�`֔>�����6HwQ�Nv ���B�/��A��u�,Ä�Cl���I�JKnah����<4ل"$��G�*���%0}�����K��[��{�_T�׿�����8�b$��f���K��� �y-Dy�9��Jx�;ߎ4s� ���(������}�9���'��R�Yڮ���UId���j:nÙ�[;�[��E,t�l��ULt�ƉNt�qx�A�7q����R�yqDD���ҀJ���q :��r���o�`��X��k���̚%'�b��!R<�F�"ȯ#T�d� ����q�)�0X k�=�%2�h2�g��7��+4�(NްQ�_ݶ����Q�_QT\��& �-���=�ܐ�GgN�#I�.ה����H�9�cN�L�>x�%|�#.�p�5�a(�u�j,Y0K�u-���[X�4}���q�]�X��V$�ta�e���_��u���-�u�5�u`�;�n��!� ��t����C��Q�<*�/�c� �v�����1P�쀋DJgm�j4�H#v��hG��u�����IԼ<^�3��z�E��J:��C�I�Q�r=�l��3 !C%r\vD��b�+{�x�3�!��,<�+�S��.�����ypy��򪫮d���!.3T1h'���A���L�1m�CJ�#Ψr�'����6,R^�j(�xH:|Fv$E/� � ^��X�`*��]ѹN���a(��Z%ء&`�{ ׵�5���xǹ�p���1�@��I�Z��(�ń	��B`ӿ���ÿ��7=�J+'�i$F��C���� �t�ηo�yWb�@T���xq/P
Bƛ��H�1_�j���{?�G�7щ�������e�̠�x��\���W��U���9���(�v��B��&�
.o_��gL�\7`�lx��Zغ��zn'��M2b"!���I�� IyE=���#�=-DM��q��S�ڧR�zeL�V��E}f�|�)�m��5�1��|����k������ ��+�h5�$ߟ�� b�]VL�h�G�����TP�����s�s� Y��V]Ƒ�"G\Orv�E��ۧ1�d'�N�&W�)^���h.C��%#.iThC����\��!�Ч7j�K!���X����<gv��A72��|�;13�"R�x-�,��10JF]�Q̞^��#X�"��vfM���Ho�˯fa]�)�jۼz�
r���꾘��`t�$�L�ص��J�7��:��c���!�Ue�ul���xJ�H��b�%@�[��1�Q�_3���ZSP�q}/��4�:#��Ư�$��L}Y1nd�*?�����40c�0�M��U�y�S�*4倅i״L$�pؽ���z�s���܂g�ۂͻ��|� ��F���t&+}����Q�/k�k@���Rx�*{<y�M������ۺT�9=���ɭ��M�6���@5��2�a�����d�a��"{�Ff4�,�ëN"���ӗ��3�X�G���rdp��T?m�ph�����M/���J�ØCQ���4�u�0jvSчM�9ِt$E��Q���fR�Y�&�۝��gZb�}T���,#)��X�1��w���g�1��� מ#M����c�fNw�n+R����?�߿�!����DNyN}�3�SV�}�j��zH�¬["ʺ�~�\�o1V��_�4D��MY�͵�{�e���~�nX�1�i��7do��z�Jy)s6{�U�Y)�eL;����#{ �b|�S���w�������\A�4��&��K&�6&J̆�sTrH�#A Y��#lֹ:����FLQ�1�i-���
L#Z��X2c���cF���[EN�WP��"�5s����܇.Ǉ.;��SsĆ�E:&�t�#0}?�����7-��_w-.:w5��?�a'���x\$d}�����Hi��}6��qe�1fӷD��"�xs~�y�xP�ǲ���h��V���R�M��W���xc_1�5�ᤓG����y���A����&j-|��[1o�\y��ȥ�¢�Ǎ?�d�����uH��z����?n�d���))�Lݡ�bNC�;��ITw����+���z�`�,��'qɹK0�A�Q1�`JX�B]�.�Ve���y�$~���xa�Q8�"�N�3>ӈ�)y%���� ��5n�U��8њ�w���"L63��,���r�u�&�	������|+�v�:���a�e�����ko�[�D��I6��zؾ� ������Y
I���JQ�q4<���T7�
<3Q>_�|���
�zH�Z�Jp*G0} ��'/ƜS��i��0V�X�����s��ǟ�w~r'�k"H���Q� .%�W�)͌^א���Kt����˞d�}	2m�4KHt�H��1#��)+��W���*��k3Fg�(��4B4��w�ͷm��c>v���("�)���)<�i2���׍y`���ų��i��t��ܖ  �D2�C!�)3#��䩒O�0.��N���a'����4�54&+2_��f����4��܄RY]�V����4�C`껚���/
cd�pȒ҈� �.���W�4}�ʹњ�!ZW��S�d�1�Fڹoi@��׆�p�	���4q���K�b��8�E5��0�U\/Y �Js)������7oze�rʔ́0��s���yӒ��G/�)+�Ț�!u��'�ڦ.1[QX��S���F �_��=��+{��d$$JGc��� aOK�93K�v�/���_��]s��.J�f�xSxveX=�&�`������e��p�/�����P�B��F(b��oʚ5�t���6�z�&��'�;ofL\,.
�-L!v�	�)٬�4dhzN���)�S�Eaw����|�j�j-��Hsk����n�3���g繌|���m\���-X6/&E�-���"kHP
��p�����ƪ�>�#i9_���U�=��锕,�{a͗�x"�c֢�m�Y��_�9m5۱̖ 	#��od�"��3�mH�h��=����;�[�,ɠ�$X�j..{��X�j>f�1e�1G�,�Z��Z��>���2�f&�e���0S��#c%�z�v�9�������(U��5[h��d�i�A�#�8W��~-H"б��\�>:+k��n�+���Zf�';bR4k"��'������`dK@���{�@"pM��H'���HDβ��t�|���?g�y�_�=U�!#|�P9�1Գ2gq�mG�Ҥz�������p��B�E4U@4���j*��>��PhV�/�Cka�y!23^
bm�ce����f��zN�њ��gJ�َ��"@O;��[�Je��/c��\x.��I8�Q�;U������ރU��Đ���m��Ny툘,�9�ۍw��o��(�/���q%����(�f��H͙p�ó�2CF����Qw=��r�]��x�dzv������瑍"�A�J6�������}�g���3v����k.p�]�M��Q���w_����P��Rc�CNd��X���{q���X=�J3.J�����C���|N;i�������)��7n���(b�!�_e�yO��7�V����`Zst��$�?�)�XY'	5ir�� ��Jy���� S��qo�yQ1�N�u"g�5�TW7�o}��R�pN�l'�����|�B-�5*D�녴 �E���<�sԵ�@��sG2�	�NdӒ� ��r��y���I(	�l���p��q�1�l���×��,��{���>��n�M��%s�𙏾�8k�X��5�6�ѱ*�~$�d�3�u��Bf�x`�"5FHR���!�L&p��*6�f�q~��H�� �`�`�u�|�0��߉�Ǒ��Q���US������C��9�8�^Ͽ��\+��p��x����P(��ן�0�����V�)q����{��E�2O-�����7{�@�ᬏ�W��s�|f�$En�$�5u���#�l��pc}xa�(�z�%��}�6na�e��dZ�E�j��
���3d��a4�����X��{+B)J�N�H��6�q�z�m�,�=M��CwC�)�����[�B��Ʋ��Qr\�94����h��6��IVW�P����{}}��hL��h�kgvb�c�5�If��:�������WB��>"8}�J�����$�u��E��Ô�Ӑ�ĳ/o��w>�#� ^��Df���S�\�)97���p7��Z�v4�ܘ��H�G*B�YmZgcÉ	��j*��[02G�׹oɝQ`Y6�� �������v�w<���;��3�c)6�ق�]���:W����Y9�J���iK����3o��WQgT\y�=9���f���8Z�N�C���0m�j��g$�i��)U��ᔟ���"׶�)g&�:#KZ"�N1.f�iJ�&�(���B����t�m��T��1c�b��f*17L)�>�	������(r�>xŹ�ȻN��>nꢊ5�l�e�Oر) cI�O�8���pJN���C��5e�%l\=��b�������#�b�Vo��vTB\X;�{mT�������/!��!'#L0�Ӗ1�{���a�a���������Ug`Xf�T�g�Sׄ�2���n�Q8B�34�(5���jn��	x��Q�d�5��&�T���=􍹐��u͊�:Ĳ��0�R���4�1,"Cͦq"5r>�c�lKw��/ݛ�(���Cɧ��]���[�P�/� �u�d� O���A�r�N	o?c)>zչX4F
�,H^;SJc�[�z�?�
&�I8�"	�D�����G�>d$�ƂZT��~��ٟi^�!�J(�Zt�^��kFe@�<�j�E��2��>����ٵ?�D*�!f�V�-Ǔ谶�x2ɮ4��6��g��J>���H$����Qx��\~�M�x� �gT+ j��<:���vc˶7�g�Q8<��u4ܶ~n�fr9ē���L%���t�[�MUc��+��1�x�_�9�J+��˲;v=�64�U�uU��\+�� U#QF��r�݃G����sF���⨘�`�� N^���[��	3��(J�@CDX���F�e�%�- Jf�;��ԋx�����$�hF�*)reS5��Ht`��A���q	>#L�}VՇ�%�`�c�Ms!������vs��&d��c������Ivӌ�L��DwA�4&��h�]����!�Q�����u�,�ZVA�ݧT�E��?��Ŀ��+<��0��!��yD���ZO���H3i|�M�+��������hL��m��-��]sVYdA�6���`�k�a�pr[.�!�fP�Eg.ǿ�͟a�{���J*;�� >�����{��Efዟ�(�y��(�"��l��#�QF����n�➗�u�$j�*�	��Ě���� ���~0�x�m����?�� �hz��"b�3��&���w��۟���`/0�5���y��m��|����O`��Ċ�� �C�R�AS���0��T@Gf�xU�!Ƣ� �d&���*��x��NL͓���#c*�چ@1�J���A��U���]��##<#�$"���d!��cGp�9��7F�[`��^��Ԍb���4���K`��;�G���|��0��m�'�:_ȑ�&~~�x��P��p��D,!�u�\�1���n�m��X0FIGd�;%�n�cq��:��(�Fp�L'������բ���y���_#E!��~z?���;�s�H�Z�	,Y܏���������ƫ6\o��%��㰋�}kV.�ik����&��[��2h|=	aPTS�RR)"��Yٙ�	j~+Yn}�v��2f|�//��h5��1�E\gv�kOKв/�����9��� �v�3AI$�t��3Γ	����FT���������Pn�t�L���,"hbB��"A�N����l<	g�]�efbx0/�>,�Oc��
~�;0z���+O�D���G&0:��g��o�
��>9�Q7%�ɉ�n�۴w�3��Dɘ��Q��Hzy�i�B*�ø����ء���\l8yfNB�YIm>��b�B�x��?�G�ۊI7��Hf�F(�ⵥ1M,)���d��v�����)|x�UƧ�iqY�4T��i��"hN�����}����� 3�f�Mĸ�Q�,3%i����~lzr3�u�o��X��4 5�v�F9a����:�P� �㲌�]��j��:���J���7�6q>��Øj����{�ť̘�@�ɪt�x��5��Hyم����9v:Ȱ[��0��SדZ=38����1%;�d]�Xh���`�p��:2c����K�T�(c�f�_��Cr�9<�b�G�	-nui��
~�FL�ˢQ��u�b-niv�_4����� ��=�o��!��>�$j�&�1v�dc5��a��/ގ��F�d]A{@�<9�Г"6�Ƅ�c	�Yy_�����s;tXDg�����jX��g)�Ș6�O�p��y��'ߍ�3xdqoPy��{��|T�;���)�Î���?7�XzP֓DZ�L3�g�a:kݕ3����3+�v�9��gP��o�Vͥ�IJ�U؁6�	̧�\�6-P�3���EwW�`K�`d�q���Y&�Ø��-E7�l�9�p��~��g߅ESKJ���l�Wu� �����Mx��ͨ�%:L#c�r檩��gZ�R9��0L�4HY j�L�<�_{��O�:�&{�mކ��.�a�OY��ql�]�G}-O��j�uLLc�9x�ykq��T���9HU�d�+9�s^F1.�'��ĝ���(^߱G��}Gp�XYX�N�g��iB��%St��YL�AS"��S�"v�qhT�c���T�R�8K��[�'��o���V�ޝ2V&���� c"�#u�h��(�M���?��5����+�<�YG��D<�c��8��8u�J�ٝ>�Cь-��Փ��Ka�Σ�^��(�R����#x��[��ΣhE��XD2WD<�C�~<ۄ��!E]�ǥ���ޚ�*"��M�.а�>�ybf�����6r�E���k�d�!���d�պ"��ص�Q��W� �JOY=_����q�4��1�x����Dw��    IDAT� O�4����kl=XG�o:�(U6V����1/I���g�kփm�)�4���+{��S���̿�O��F:F��$�a�ڍcx不��?y!���a��#τǀ���ǃ�����i�W��U��?>�~����*r���߫���Y�~��~|������J�|g���k_���0SF����o)o$=�L����Ӝ�F�g���w�,�k���Seugd-@�Z����HC�Ⱦ�������2D��h�fS0�4�����s23�s��� 7���6��0�:-8�e :@ſ��k��O�,�2��<l��i�`}*rb��F��f���L1���B�?k�Ʒ��"�⹣,�4��J)o�=.��ڋW	0�V�oz~����<T���>�	c�a�.0�\��k��������g�8$�Yq�%;)�5�.M�kv�C�v���w���<%��dZ6+{�'���.��3Ob&�i"کc����ֿ�Fr����nz� ���_b��*҉$��:�G��W^z6��bJ%�'�]�}���w@w��E�y����~�n�|���;Y16�Kl��P�a���N`�m�i�l@2�ś���<�Tk3�.���+�z�:�� Sn�	1.J�G
�v�m>�;x��@��C4�/4�S4���,��[�tV$�˪�-��Tr������|E%Ԝ5���|�,�:8#PG��@>��Ջ��%X�r��N����NG�7��ݎ��KX��������16�I�3�h���.Z{�e�-��~4K�0��;*?�붮��u�E/��	��V�J(߇L�����ukV�^�S�`���L"�\����Ɠ/����y/?Z@:7$�_B�:���sA,>�Y�L�RZHZ��M��;a�*��;,���8�G+�G�1����`ޜ~��M5�23�*�!�I���"�xv���{�w��vfD�yѤ���s-0gm�q��R⧎ٺ�JG��	0,���K��t�!d
KLɘ&�ʘ�|���p�5ua����R�j��ZNK6��P?�}1?�F)����Y�h�vG����q�4�A���+0�ז�	2�:��A�T�b�ck�1ոʫ��&�R	�e����u�INܘ�S����DP7ԏ]sV.�� ���Y%������"��:u�W-G6��i'��Q��������.��*�4�A	�n��/}�r�����JC$��5���TrΉ�&7C�ܱAUk�0Ym`��1|��;�Ɓ2<�ΎId�9]��ʹ�U���G�L������,�{�ɘ:�_�U�m~�=�-���G�c)$d�A%�L���෯�;?�N{@�)�٬����d�y�5�7��A[x�ϕ1fú��y]+ULe�J
z2vV����2��ܪ��z������t
�廄Ϗ]G
t�|�V�Fa���ͦ����Z4ʽf��"�_\�׽o�G�'�J��	�ؠٺ��[�|O�i'�"�~���5���D))C*�� +S��B�\'ٯ�Ūi�^o^WsR��#p�4�&��[��I���1OPs���3ځ�P��,� �Ր��lglX�3�/�ikc�HDb�I�HF��u�9�<C��N���l��-���+�����ؽ�(��"��!+�]��N*+K�*T%�ʙ�q9T��F�(`�Y<4,8�uC7�9d���F�eU;ٽ�S5�2#FN�����ͼc��D����u�<�D
˜I3��k$��̦	,q(>ǅ�8���us�(fbX4oV.�+u�i�V`�̂���F��R���-� C����1<�؟���[���d~HFl�j�t��U�{���U!�F�n�
��uki�	�Q����[�����5�
G6�S eK-��Y�y��(Rw�@�Mt�\ѭ!���<>�f��2�.Ƨ��J�/�����#�X<� �ܻ߿�!��!�LL{��mD��dM�z^�0��]�5���xݺ-@�=�{��=�\\zޚ�6S�QI�h>�Hky�[���A΍������'�ŗ��&-��[�Z�"hU��Tq����߉��q�4xu=u/L`�~�7�� ��:�N�`��a|�?��7�A��G�"Q1?��=���ߋ�r�t?�}�FjkZ��m��9�=��S��U�M�Pn�J!����QȾ`"�d������n� SaL��L��>D9cJ�K8V�Rbʜct��Q�9�,qΘ֛2?O�͏�2h�S�1,�}Ҙ0���j4�4h�� 1�I#�K�����c�e*i��D�}�1���Y@	���$r����.õ�7�i1�Θnɘ:-�X8�����S�1偷�P����x���{1��yd�Y��R���.�|�ϴ}xn��t������%CQ"ĉ�a���G:W@2�s8��r�]��1:.:^	��<����S��q���g៾}7�6�I%ql� �֜� ���/�����2¢����q�������9{>r��X�t
��q�v��80�@��c��~#/$�]x��nbک�X\�ZD�qP�H��/^w�Ρ��zj�,�CI�(D�b�R�"������eT�,��A����)5>"ؓ�Y��PJ!�B���
㠦��D�jK�N���C���.����8$;.2qO���Y�X�|!N߰s�0�HbQxX�M:��~����a���Pj�p�XG�]4[|����JX�H����KTqԲ �fzk@��%���i�A�8�b1W�~�]E�t���k����l��&��
��LAB��(;>���#��wOa˼f��AB^+�{�t:&���!oc�fJ�M!,�(�3)u<�!h;%��	$��8{�l|�������@�Y���J�Hcƈp�5J�k?�:�{�&�9����y�);���J�Y�?�2`Ås,�ENf���guv�la9�&C��3�vL�Hr�f	�	(�V�V)�����T������$0�KÞ8�aL%4h#C���r��p��|kf��T\��@�ke�C%���錩KWަ'��2�F%�ύv���o��	��f�4��h���*���Kp�i'a�aL�2 N۶����^߼cccR�L�5_v1֬;����݇ߍM���H4��"�ɉ��x�.8u!���waƀ��1�X����Ͽ���u�+n_��=���c���'��D�F���+sޯlُ�O��@0_� %%̾�!�K#����,��CS���?o֯�%�/3{�V�5TZ����K��NF0PH���nf�y�O�|7�r/����l�y�v�mA�+�w�6P�Y�]���њ��7�g��2�����ݦ����,O(�4F�ica��m�"�5��5lc�C�U����ḡ�Q���1��o"�2>��S�נȳ��1��k$A����$~t�}xy�Q4ڔ���W3t�W��V���D�ڰ��e-��e^�NU.�[×�Rh[�vQ�4r�Ջ�x��^�5KQ��d��bB��-T+��E��Is���7�u�1<��+5�<�?���J��;��8��k;�����]{���(&�MxT�$(/O!�H�C�A6��Y).�ܰF	%'��2/M?�9+�=ja9�1�eE���="���G.߻���i[H֜���&7��(�6 ,زŵJō>4���b�?W+դC��%�\!c-�t.k<�w���F�H�3��Y��;���k�RU��`*,�i�[/�U�����x���x�[�}�qԽ4��3D=D)����(�k(�ԣZ�K��4�����R�:��Vf�$dC�&e�	mA�����w�8�����S�XCȚ4{���xO���T�U�,�!ꗰtN?>r�;p��֠�3 ���O@��������fk$�b��m�Y5G�����Q�tE݆����AUw8� 볇g��Ѻo�5�i,���r�*���i��V��{�5���;C��ݍ���|�+���P��Qi0m��v}��!��ߏ/�յ����HQ	A��\n���p���x߿�v:4��W/�?�ظ~6�R�I,$��n�Ov����1e��G��Q�K��Խt�2�>O�/u�]t���B�.�>�'*A�����
��v�4��xf;.�J-��,��TQ���(Ee�}��0��?���4OL�tМ,��pt�4�W�H!�R�XD�du�׽F��<�(bT��"��dFո�fy� a��t�Fd�4bU��2��2�����$>�Kpͅ+�όi��w��'0��ևq����|,�?���{q���w`��߃z����!�NA��Q.ѮG�q�">�*`ddX�FnȌG��j��,�\k����8��� �M��0�6�7/h���k���8�Y���~ZS�m����߾�;9�/�Ş�[Ѩ�!��`�pkW/�[�X���������Wv��]�mRSF�����144����:^�~��>7H!�-����.��չ��-�|Rx�!��}��Vc�N�X�G���u���AZ��w�4�n���
���"x��C��ïH�jEq���Y�$[��R1�:��M��g�qN�ez����*��y8th��@:�B.�<f�c�X�r1�OF:E��v�÷o�1��\,Z�7���U>�D�ّ�=!$s���I��*�B�@R�v��9��*�aB�4�B
�b�M�:�1Jfh�%��Gџn���mę��A_>��sg���=��i妏�<�$��)�k0-�B��yǨDx��%���j9���R	�};r�(Sɱ0Ƥ�x�`�nO"R{g���k�<����p��7ҍ
�:�[+�i$�v��G�݁��ql?�"�7�gL���+J��^*f6�Aa���9u��y����4kZ�~�q�Ɗ�S�	
�<�-^����ru�Kĕ�9�E�0��.Y�pƌ���);���T��jux͖ܓ�@�)E�3	x���#�ꌋ����bmn�m��*���O`�Nv���4�0�I�y�@r�?k�SC�YF�z�vӆ�ҟE_!�J����
�=�Z�*�,�.&�r�2c�X���)h�1��uX�T���h����:@��~�|�c�
0���Hy���{�y�9s�Z���غu;{�	8xD�)��BS������A��ct��J�!�T��s%xOLk׮Ɔ�'��(a��ر}3J�1���D׾�J|�C�G6�ξa�l���ֽ�����t12�Ç�%f�L/9��p˯^�܇f����4)2!�k����>��e�?���u�a\{��� 1.��.[`�;O*N��{k�ΒYv�_'��4{��/{�i`Y9��|��ʷ����)5g���0�@IxOhP��'p��a|���T��F�����~�l�WA�G$Q��H6�xp|E2c-3$�'>l�)X�5�1�k]o�a-<�u��0�F� o�ʕ��x��O�E������
��WJǭ�sk܊����N[�W]v>֮Ɛ��[���s��-�(6�;@�	>VǶ������/mC���o3�0/��`��J.6�0Ṫ9�ZXZ�Y�Mm�J#P�}M�0�V�ĢA�Ѻ�Z?:�[��w���JI�,�*�z�����i�=}��W�g#�js?Ġ����|�BWZ3߫�>:����
�}�A���ӏj$�Y�S�h�V�d����õW_��'-��)9��k�)�6՞�r.�TQ�z�����.<�ċؽ���Z[#��fι^Fd���2V�RȤt(O5�*���|ژ��i+�h�F�X�5EC]�h=:�2k�i���i��hMFl���g�M1DՉ�R�d\u�y��5�a�(ex}X�Pi��k���[Q�2�mjơdt��o�-X�WHmdv$݄�$��.���\H	3����5B��φ�!W�r�r�u�Ze|��⺫N�����R�A��~�"~��?���D�D��x�Qx�p��º�����A��q�̍[�8_�]+�U���?���X8�������"#���( ~��������X%*�4�7�T6+y��%Yݞg��waS��K��,<Ox��������j=Ƴ-���U�&t;���2���h7�0O�b�6|��Wޔ�@���l�d�k�L"�Z�q��1`IƳ�C'����Z��R^>b~$�5@��FSL�ZlZ�ˤ���ĒI1̲�BHک8��,B���Z��x�;�c��4c�u(䈀q1?��&��ߡ��|�T|�S�9���A���ރ�^��b��t4�V�&YL����4f���5K�`�tL�6�)S��(�#��B���	��w/mލ�^{�5�Ï���ɚ��'�J��U��D+`t��X?���Ob�̘rN���G��ñIO�����
&�B�S�A�L�UW���]�6Tp)��u��M����5��=���'_A١v /�Zaxy�0�@�5t֊]0�^a!���<DE�@�%h�QLH;X�h��k1Td�k��z�14r�V4
�k㍃���S[��q�<T�D��H���)a��v�A�L���v�s �q�%�ν|�23���f��c�f��4h�/���\ғ�h.E6�@##CD��;v�'�����\�:��&��Qs;�ē"���-b�8ē	$3V�@��7QΥ��݀�4�$�E��s����I�8�*����vp��o��u�PȦ084����ƟD��8�{�Y�꾧�mϘlR���Ĕ����b@�L,�x�	f�Y�����(�*%�-��DdC̔�<�i��T{��8k�l����aެ"����I+3)o�)�=yt"y<��v���Ǳ�d�<�6l����H$�d\U��3j�d*_9r�������5��u�.�J���Q�b1��P�J}�1R`JF[�bL�
Z�+q ��>D��%���y�\J��'�m�Y�i��@�Z��t����}H��7�]�hD�)YS�s�p����]`*Rpn�Ʉ�`����+Ɂm�3�,�m�<��f��8|�Qb�́�(�\&��$3x�`���:pZ�kwRI�Gd^���K��o*��(O�(��H�S�q�9+���^��@Q9�2q��*��<R잚����2�q�`��C�����ǒ�1g�,�u��q ۶���D�l}}���j�*���b�s:N?c�})�k5l޶�o݊׷n��۶�3N�W���K�E���2tE^�q�r�-���`��~����y)^�9%���K��OD#�#�,�+"��D�!�Ok��L'��1�a���ghb���� +cb�' *�;C�^Ȧ
�ӛh�D�@0-�4��N��
q��M��{�{����fKKQ�5�Sq��0%��=��������%�ؒ}����������ᵓH��K�Q��-ňy�tDB�{�eK-`2/4U1\��0�`�Hq����try�\����K×{@�E�ـ��&�F��=̞��y��ۀSN��)��05c9�%a�4C�ҦO#;�ş^݉���¾�c�;�D)1N+c|�*�8��Ld�LeB�����iE5���o�Y�e�U��[]� %�Fr]�JAufRҜ��Wx6��`�kGW�����C��Rs��B %��J���y�
��rki��}aH��d�F~/1$��/I����qD��Qs���sO�٧����`d �,�5��0`F�,��(4�CX�2�������Җ��3p��,qDSI�CN0|�;��RVKbt�bH����FF(��e�e�Ԛp�<i����j�z<:��Z�����8bm�	�]$J�F��1��QdbM�{�j\}��X4o:
y�^���q��O���Ӧ���z��Pv�Af���`��(�Np��q�Q]Q�_Y���K�hc�d?3 4�hw]kcq�R8p�5����2>��+����C��Ö��/�����e��Ы�he��r�cI�
Q���(܆hs�M��|����̥*�5`�fO�N�����U����r�<$c
��������w�X-�Xv����P~���@?Y#���1y��]����D�-�v������	�g����`���'�+��a�C�y��sGfC=�����4RȠ����������`Z�`*�D1�A�������U}�@�Ӗ�1���3.�^W`+�7��guJ    IDAT��+1���֪���6�b:����-�/R�g>p)���N�L��w܇�는��� �^K`ꡉv��ݏGy^#@.���M���Q�~�*\r�yX�v)�OK!�f��韸��E��
��潸w���s�Q���@�&C)�g��z���WE�]�,�׿�I��=F�~�Hy���Pȥ�c�khV��Qv��y��Kp���`��	�n�1Թ(�^����&��_a�1 QD��ns�dj���y�NY|�mK��4�4��RzXC�6��BÅ6��Ŀ~�(2�I���L'Ƹ�h�(m�� �l?��{'���x�`%�:dm.\��E����5�����
����?�ZT5�2Hzi�Lۧ3����L���1�.`��@�L�|��j��D�k�f�Iy�����s�d�t�Y��82�֊��U�T��l����s}��!������~���˘K�Wl��3Ev����8u8N�T#Sr�G��q�#xߕ��܍P,��L"�J�d�T�aǾ�x��?�����x�Ga`��30Y	Pm�(���5�0�r�*�������� g� w�H��V�~J�<D�:��8�&K8s�\���31gF�}gY���P`�BIrc9����v�t���1��$go(����x�0�'H%2F��F�i�8Ao��E�r�a��v�i8�(��f�U_�]yd��a_�y�9[��z�c*�.2�,���	���Z愬q����3��G�ͺ���2�}H`jS/b`���vb:l��$u�� �)�g�y	S�c#J���<l�q�6�Q�8��G����"�y	�d�1�tz�r�1of/^�ta �Fo���&�qΓ뛊�ր�\|�*|��bjQ�pU1X9�)����]/����,F�NG*�B!��3��z��=;��*"��"��ʳ�1	vEitB�������H�c�b���:ؽ����K�3{�=�1s
%n~��t��*����$�q��~|��>���R��9I�_��� �<�y�b����h����)��_ׯ���fR�dw����r�K쑘3�J�1'�L�����&3Rq��IU�OA����N�vS�F�u�?�P*�z'�[�����kץp]4�sg#�M�Vwp��8��@<;U��Z��c����?�]�-���"0ձ�M܄u�L� 2"`���t-dW���=�{���;)�y�L:�\qڭ��S+�Y�D$�a�p����,�Z2�)E�,O]k.24��[)(�Uؼ�0^xm�l?�����q�b^0M��H� �A�J�QG]�GV���x%!�{8us�¿�1	s��O�j+��� �'�&�͹�s̞�Ë�77zF;��}6���K����Tי�+m3F�Ϭ)�]�v����&�� O��Eٰ�Z�ugP�f�FE���&�L�a��E8y�<�[�+���`3��)�1�	�cϽ��B��=��MO����~{��(�,I��4��"�ec�J;�1�J�-�2̠y"O��o޽a�������Y��K�6���*�*q�k%� U^�JE���/3ԍ�8Z�I��:f�`�9�24$�g��Q�:�@3`Ӊ��o����Ci�ۆ��Q�I�9�C�cW1kWֵ���1�����$�(7�����8��ߓ0��Jy��*>�w��� 1!V����������~�<j(�O�	0M����jp&��q|?�8�X3��ጵ�Ŭ���G���nڕZ�}idӤ2��k�"R�{cZ�0�+o<�V^Q�9�U6����Ɯ�&R}�]Ky=�J�OL��� G��=��/s�62�~��T��y�h>��BQ��%)6�V����tO�K�����qQ;>���+�̘`JƔD����S�� )6����Θ�<�b~�Ӹƪ�}Q�e��9(�v���a]D���^��_��ǘ����n�������\2�����Li��ރ�~~�G����x���7�����j�[36��m�m!�E��!�E��?�ĝ�}�nz��9yʀY���Σ<n眾������O�0��~��-1�9�Юb�p�����+�&n}��-�[����:��:���l�7	?�C�]�_�Jeu�TA� T�R����lg|t��h����|��q�i+���ʫ<L�M���LĄ��!�vD,�_�v���ع�ju��I�0�Kɧ$��5Y@��\d
C2s(_�EBu%���9�I���14J�HD|�#R�6�/��%g �$8�LIK~n��L;�,���-0c�L�_��t?��<��n�=R����P�<.s�����g�I�o��h1�<�VP�"��Y#m��N�Ӏ�j�4~D��ՑI�18��@_�V	�����c� ��J�hy.���&�&�80:7�\Q��.��u����v�C$��"�V-�R)�9<��b� �S�1�	Jƃ��p1q���1;p�F�
�*Ҥ8m�t\qљ8e�Rd��0�2b�׭�FL�t�5hGq�pw���G�-��cE���>��4`N��j��8�,�iF��jX-�9<S�[��p�2.��L�k�fkш���m9��@5�eLi?N��m:He���ˁo�qTl��Z�:��CG_f�����)͏�I�zH�!9ҏN6)?�y_�l%x����^$#	D[�Hy۔�ҁ�2an���(h��{��K�w�[U][�����R슊��{C5E�)��彔�DM�iv��$��@�b�����{��1�Z��k����$|*�{�9{���s�b���Q;�^R��n�Q���E��1�=4W9�T��/�Ǎ��F�ٰ��),��p8�Q�Gb䘑p���z�ݭx}�j����*��|��L��{p��S��ĐF�mJ~�9)�>F�s��>��ׇ��&i�)�3�A��ѲB���i���uZx�4���5i6g��)��� ����qgw�>���j��!����/���ap�}�dTS���.E�ؤ��E��I"ň>���'F/
�n��a�~P�q�\�o��r�*L턤FS�M�����ŉ� �>º��'i���]�8[*�_�=?;n�y#���+Y`m+G�;�ht%�ڕ��,|�[(�e��>��xBҠ�iJrj�k�-��#�M�E��24�~q1�:��E���kg���/�3��?_�	�^��V�ȥR�\�&�P-���p�QS1紙8dھ�"f�}�R-��יE'c��Y`��N���2|�|���Q({� .�����4�'N��N�c3%���#��kij��P�f5�u��,�zz�3!u�ӺW:�X"D�����ę�:{�C�4k��["s����sk��FJH]�#�b��1�՗�nT�:�&i�u�X���ȟ�L�ƌr��@���\6)�J�@%-��Nߊ�����=��Z�g5�}�<��D��ƈ��5��V�aޢ�0��Зv��m@��O��9��y�.��E�h�F�iiKցjΓ��i�����-�>�}E��U�,�R0�tM��#��΄�"H�T\j:���{"l��4���Eɿ5Xv���p8�v��Z��k�.���_�v|�>��[~m�j�2���P�����$0-��rep���𝳦�׌dd�$��c/ӌh>ҮT-ȑ	�`ö�r>�|���.��9c����p������T�q�ֵ�n{�*v��јrb*T^L#�-��T�*�E�6˹�5�����3ԍ�<��mW*��9���	�P�n#���43X�T%�Kjn��Bi�H���! =y"@CURֽ*+S�i(�M� "��2YLsJ�%��Q&��W�(�+砭J[1H}�ߢ1ͤ��yF`�g`�@-��2��1�����Z����T���^�n���=I���b�<}H�-�<p�/�/�)��F���/���F�d-9�n��o�Ûo~�J�W!���G�����\�U�nQrÌ��)X�c�S�өn4O<��~�]�l�K�d�DØ�$���Q-�������B�RӜi�N�r��ؾ'�D<�d��P	�>���%2y���r�8��5��Ŗr1>0����4"-c��RǠ@Os��ZEW?)�����ɘ�ja��6�D<�!��E���Y�]s�dk�^z��g�P�	�Wn؉�?[��[��ig��<�	�$�8p�xL��/�~�9l�ú�	$�l-S'��3��G�\yn%�^:�BZL��yw�8L7R� �\6b��lc������ԉ)A�5	�um��nu<\�.��?��\�ٲ��������E$��n��^lۛFg���7"FX<<�<\���'k���*��h
V�s���2��C��A_�.�ӝh��᧱L6�L&m���34�p��G�c���?�|�t�Z"n2Y:A�1��Qr[���欅Qv����qK�]B��Yu��F���h�b�O�][\8���q�Eg`�6�IH�~���
q-�t�_FK�܅�lƢ�7bWWْ���7r�Yv��@0��� �?$��M7��!���+��Xu2t�uB���Q:-͏*4)3��Ǒ��-����������*6W��*I�VN����狨��Bj	'��7��	 R�ZZ��թU���V�����&PMe��W����T3����k�m
'����3i�ݒ�#��~s6���'h�^�R�l��J�so� x���~h�R^�%Y�rN\Ǒ������\}QG'���6���KE�N:�D*��С�E��OK�g�c&���?G��:��/�%YS8q��4f����3r�,Zژ�K%]�� �=V�폼���a�&��!�W�����C�|!�4U� �0 M-�x�	��q�����`�b*G��'#I0n�l@z�Q�㜫��N���Q+�j{�)RL�o���*���V�6�P�����K�����PC���R�����S-��"x�\Eu�+��(��ō]�%��i�>P����5?_��qh7Y	�7L���"׃J�3	��n�|��,5�iR9��g��I+�Q-�7]�3(1�ݗǌ)cqť�q�64=��n�B�<K�a+��F%#y|��:�[��w �w��o �a�5 �g��e7����^��k�I��qx�N�j~�}t����gLcs�����i6�^(���0�O-�4OLkM"ۈr��������������sG:�N5�S>�y����լ���(ar�����������4fV6vE< ��S�[�U1�@>�#gb�]���G�Sg�#�c��4�7�]��� �|�4/_hS�b}O��}�\��/]lBp��G�M5�z�Y��m.��jt��ّ�� ��.��vM�ǧ�.��pM7�ڳc�&�ؙ!yl���9,>V
�H%�I�Or�i���/,8�� Ӻ�w;mw2��n��YQ����-V��+��_�8r�.�c����S6{i��)p��B���U�����V`Zk�*Cqɚ"��՝�+4��d��PS*nz����GƟt�����s>`���
�H34����rM��T���������D��Qt���aV˺�\^O�Y�o՚kd�dj��69�&�M�bH������ԋ>�"^��*(��f��gK������0*��v�d(�t�#�J��� 0�f���F%����n����G%��Q)��݌�KDЪ��2�2J��L���-'��<�]P��V�>��dMScڀ>����p�1?��A��f���јv�[�{���H@�I�q�Usq���*�{q������?��Lk�2�����6}���iW�ҭj�m���-G�} 5�:�1k��>�s�|�ξ���P�B� �^dr	�*}8�؉L�Ĕ�OV���;_��-�H���gz1fd#~���`ά�c���U�cwz���
�΢|��cF`��Vd|��6d�@O*��"�Q޸y�E{Ƈ�R�0s��؅l�߹�,\q�hk��/�c��ؽs�踆n��V��}�z���]�x�:,xoVm������U̥�����U�⨃���S���
���a͖^�]4�"ȿ��[Nߕm�W��B�-�"��u�q�4�M��$+����p��H8�YZ��=D\rplٕ�c�.��w�Jj6Ǒ��k�}F�k��3�{w�����N{n(	7%%,�$/Ul�S�W38���p�	�`���H'�شiV�X�ޞ�Ն}F�@��B(M`S*!_, ��őˍp0�}���&LF��3/�潇d�*΃G2�Z�̨+#W�`��x�ݕ�IІ�Zv��pQ���PY���\�?>��Ѿ�7���}��3���Ǐ֘�y�S�8�"�ocAlڑ���Ƈk����IfX0P�~����q#�����+WoG<�B(�@B��Om�dY�&���3��HI�,f�1�3.����pji�l�f�)���L��|� �Z�m
��^:p�&L����uc+�`J*�l�lJ���6"`͏��U�TF���H�5��n�sb����	0e4ZX�����{�S{|��и�|�aO����y�pD��c��z۵H�z_�1���e!�s�kǝ-D�Ԉ|�^U����pʬ)��;�JCMuOЃ�5em�	&׬Y#T�	'
�ӂ�1+.ɁMtuK�s����m��T���I�2)٣Im�G5*��ݺ��хϗ.����D�(��-�rWo	�?�V�ـ�#[q�w�b�Ш�ܷz3���.�O.B�F�a �����\��A�TD�TthBZ�j�����I�ɿ���d�
�,f��sʹ��?�:���hE�O��]�G���_���r�#��]f�,q	���=t��g�Z��uҢ��m
T�D��X�Т�L�FN�t�1q1��˩a�Xɉ���t���6Z�����
�q��~vU_Bh�j''_�v�:��L��j��B&�|��l/��<�8'Μ�f��C=RO������w����d���M1�\�K��Ǫ�;�ϣXe��))��,Y	D%���23-���4]�+���=��z���m��ґ�ic���\B)m�4ĺn;���1�]������T 2}�5L*�Y׵f�������L��"�M�/���j���d�.���:P%	~�i5���Vj�V��6b�~$,2q�W�7/������U�-3�M|��J�8��"���9d
�>d2���(#�LM$����Ԛ�0N�'	���,x�s|�b:b%�}p��F����+����$��P�f'`�qT�S���Y�3���6�SۨQF�JEd�2��12���g����H�x��	�� łm����DہfNmQkW����YR]v"\�QԭC#q���q���r.�J������es��.:m���7�g���1B�x����HP���f�KR<���!S����ԇç��U�<�4aC�W��9l����k����|���E��!���0-�=V�+52��}��X,8�<�`t����?/(ഔFtB��0^�'�6�2��4�P�����3�F�~x�t��%ZjeQ���%S.4�z}��O�����#�/�Q����%3ްw�=C>Nni6IFMm�)a�1���S6�$��0䌉�=�-0%��I9D)o1�W��{
.���b
�*Ƀ������z��h0�}�q�PYDi _���]����,����~���o��SO8L�֔hu_9��A�pZ�Fj:nR�S^�n���拖��o�%�4iny1��׏��?��]4*/A��}��]/b��)dS]�v�p����p؄&�קH���[p���bպ-b�$YA��N?�k����E[�'��]����w�ݜB�� ��X<�)�c���Xj�J�voY�j�7��{���C4�R1_F{{֮Y�I�ø}F��(MQb$�.|�<��'k���vbö�ک/�q�����q5&�m�b�[��]%�����t���a��N9e@��<>�/1H���|r/Ə
ᆟ_��c|�/>k��c(
5b�C��s����&���V$;�h�vvT��?�ͷ�������9G��K�C���8�i��;Kzq�#�iOF��H    IDAT�H<~~N��n���qZ��џ�����gOCsH]�����ġ��uc�}�������:Ҫݵ�����ž4���?�c�-@���rW�=߹�1k��@�O����.Ď�9��Ԃ���ݾG4��=g��`� ���>}"A��+�7��G!���#���+�������PCL�<ز3�����[������>c<�>c�N$+io7����X��*�QwI*.ؙ+2SX�Y)ǥ 6Sua�ߤ�zF	�����F�xPc�-��S���,6���3���l<�l&#���.�Y�M攗�&�ĸ��W&��� <@ÿy����`JPjmBh`�Ac~�hv��a�Z��7Aeť9�1�^��
5_�+��d(q,�hQP@`J�
f4�6�����p��mh0�������Lcf�Q^� ���=����(��,�P,fદQ��0��5�a@C�����E��D�|�)ZZ[1}�tSHk�K]�]�ݾɎND����Di�e�LJH�v"�N�[k0��a#�4�&G:�vb��y�y�L��o�t�x�����"n}�|�b5&���^{9���·GUw���s��V�F"m�)j��<���)W#i�`�)��Y��Uhy�B�?�˙tI��&���|��u�-�̒娟���� ]ډ�0�,'
�F�׫g�n\�w�-�Dcm�Au�eET"�щ���J)�L[��~v-�HU���	8�^j�:h��^�yS�i��([��yP�����dI��f9�;[��aWHw�1T�)�f��9�0~tM!e�YM�\��{��p�$>X�|�[wv#S�&�َ�+N���GW�7�	p	j��i������ko��u47%�>u�\j=y�M�gr�%������T&Ԃ5��#���i�#V�(�!?�}�M�SK�Jp�2�F��d�GP�q ����B�c'�U��SK�����JX�}Ln���(��4Zd$R!�R!�J>�`5�Q�pܡࢳOƤ���?�,�)ݫMk�5���uOo�?1O�%O�x]�!�-�a�4'4>I���ëo�:,1a�a�ר�i���֙�6m�6�~d#M�:Vyvm�Y4��*� 3y7�N�
p�3l�����ɹuְ�[�\���i�|.�õ�3�c�5�,��X�gnu��|I�4m+�(���WIc�������`�|+�Z� xn���r�,�x#��A�!,T6��0��.�R�\鞝�f;0}�0���k1i\3�L�0Mb-All�N�yw	L}i-n}�etg4B � `Or���ƃ���N�6X3ى���+�ݘ��G�	B���s�q1!�����Ԛ��t�\&���l�4'�Ym:s�И-�;B��Z�f\qY_PF���Ĕ����F�P�vd�F�*S��Ք�N����U*[�<UzydRIm>QH'L�s#�)��l���x��i��4�H�߿�T|���%ǴX�V	�H���������>y���:i��vH=�bu7��Y|����I\z�)���a��PE��Uh���mGǩ�:ٲߘ�&�gѶ
?�@(�E�C�s��&+TޓgM�-7|d��Tc�|c7��<V�ݍ,�l�N}�~��o�F����^,[�7��a,�b=���L�*���2f�>������M}��}��������Ѽf�j3�9D�>ʉi���7�A9Չ?�p=�y����K:���ưp�"0 �?K���{w��B��_��o}�k7w`Ն��Md�L%Q��pȴ1��?���������yx���(��B�j� !Y|j�R(Ĥ�UΣ�jǡS�7?�6�v������k�
ux��c����g1Sۻ.��H��g���ے����O��:i(Pg�K/�)C�9|�L���>��۳p�[��c�yh�c��j߉��������}&�9m�tU�֕����-�-hi
��Im2�/�n1�� ��[�ߟy/������{���{���C�rO$�����q��o`gw	�jP&Ӂ�O4�E	�,�N����������Ł��3�y��g˱z�hk�	��� ��κ��8.q�]�f�/��fc�z�Y|�b�E`��p�5b����trǉ¦]�]���ݝ%�Hqr{EgHZs�9U��M�蚕�P+��5'8L	F}tS�PfcB�K5Q�8�	���t�4���D[��f�Y�fZʃA&�"E�Z�����2t;��5K*oS#B�Q�Q䴏`�T^jLő�%z_������Q��t]�	�������Z��m9[�쪢HjL�M�2N�5�>�Ct.6�EtP��e����Pm�oq�O���>�>|�a(0-"_L4?���������j;��W��=x��w0r�(~��vL`B��ޭ�۱��&Z��]�%ϖ�]��� e�m#� �:PM� ܾm^z�E��g,��y4j�|H���.�,d��5�4~0~x��7�Q��@����X��X�l��Hᨸj'��pӤ�g�L'̔��"'�
"X�7�<d��S;�v����"i���Ӛ�hS7�Km'�z���mrg�Z?�U�RG��Oc���_��|��>k��:`�c�:�JIje&sR'��I���9�;kAiH�7`��Ψ��Ə�W`-�"alSD&XVz����f#�8t�M����9T�����Y�y�>h�:����5W�6<��p�M�]�e���|�d5���E���O5���s�#�ܙ��U4S,�pY��ՃR��QgZ@Skh�5b�����L���������F3�!b������L�I� �����Yh33�۩�D�������m���sV�N�`e���g��'1o��X��/5w�Y�NXE�g�y��1K��r>�r���q��)�ڌ٧�ӿ~Ǝ#j&n�!�Gߵm��$=��Ӈ�\���lB����2AAm��TM"���!8��:�ם�>sC�9?k:_�а��^3eN��h�k1+z�u�/�K���[�ۜޜ����w0�)�]/�Fm��c�����A;���պ���0�Sw�$m�
Ly*���F��ǨV/~���p��(��B���s�C�M��x�EX��6d\-��^(���ަ�!���܅x�6 �%L��4q��`2;��-�|���G_\��~=y?|�6	K�;�Yզ$#ڸ`SE��Lc�L�6����A��w0(��1�'�J�W���hb��\N$7t&��c��>����
L>�[�uj9�dy�6��L��a�i^���F��s�Y�&�S�I.\��j�j1�E:���9�ʅa��U\yͳ�[=?��)I)��%�r�r�R7��{2�y��t+w�_�`Z�|�U<��")�O��\})fL"Q�,��w��$>��c�*��o���8�1%�Mw,a�v���O�7$`����I���g�ٗ{�+��Kf��Q/@��N=qn�͕�Y��.�ǯ�����-�T��8x<~�˫q�>!�-�;Uo�����'硷��PM
5�?��%�����������O`���	]|@ęU�L�()��M`�i��ݸ���+.>~�A� ���i��(+8�c��1b�$�?ӥΓjZ(!��b��.,_�	�u�;V@W,���t�v����੣����M*�1�=}�Mw��;�nF�#��4�&h��g� �/�&I�͢�ً��G�W�_�1m.���)�Wo���0��Y�aZ[�[l��xఀ���:{ e�
U���˵;���/�y[��*�6zp��Gb��	H��c _u��/�p�Oc��4\�� ��!Ɉ�=��ڋ�=;�)f1�Ʌ_5�9X��i4D���c����6cG�I�jC�~��n�\{���ʝx�����G˱���`?��E���S�)�"��Ow���cO�K)C���r�qrW�K�^�g;&���W?��'�A�{;z�`�������N8�'폀_ו�I��O�@Kl۱�wv#���p�"z�	4u<���L
6A�y���v�����nx��2I,�s��M&mch��A6�9o7����+�SS���
��S�e���L�DL~f ���W���@,�s.N�IF�pjZ�.�'�7��.qѥ�[��,�%�)� �4@R�j��N^UdLI�5�@�^�<x��C]�d�ʶ�ϸq���،�8W)	���C���O�x-Kq��r��у��=����$����Y��e/�x���d�Nx|-�x��dR(P�\N�����'��:�Qk�b��Y?`�Bgg7�y�}<3g΄׫�C�ܟ�%t�ۀlG� SO8���BA���PЇB.%Y����%4�p� ���T��m[��g��kv�'a�S����'��*���<�X���ӊk�<c�4���1�AO���%x��Ȼ�#<�6ag�!�FϦ�,�i`��Z�=�PUPa�
���LA�Ы/��6�GM'Z�XS����	��>���b'���Z���S��ø0�瀚ﵓT���a�u�5�Ѳi	f$5fsSF�v��t�6�+�|v���y�_�5;�G]ca�$��.L�=��RQ���d/J�^4�*8m�\8g&��6瀁��	U�*%15*��s���xm��ض'�tɋ��u�e\�4�H;��:���ZJ��ܚ�Xg~�Z9y�9{�]K��0�pu�5q9�Y9�S���Ȝ��{b���7\G���J�4�|q�1�:��&�ș���6'�n�>bIl��T;z��4cL���k��FO+k�\J}o�2sc �\8l���_&S�F���c�s���<���u\1�tw�k�	uS�J���Gc�x�yF��^~s�|e1���b�60���u�Q�UӜt�k�[��F�R���S"c�s�����1�S��D��޾���{�H��)�����@ߋ2�4K�h �M�e����>e����g�;K�����}���^���LJ�=�T�j*h'�U�F�@�a���!����k�b°�:��{4��p��t��n}�M,]߃��eO��Dl6�e(�){1�D�o/�}{��p�Q��:3&uh�N���Vqy�6���p�#��+i0�:�
T�����#���|����zsf��3�Y�|O:D������R`�c��ZG�i��o�U^�aҜ�����"�5UZ@`��!�8�tFdS�|�q��5DQi�@I�����Vc�o�L".S��Q:ǒW�1�~u{��3SR�����M�$�����ݸ���qř�����T�V	{J�ݏ��?�{C\H�4?��R̘8X�U�
|�l7n��q,�d	F���;�S��ǇX� _��ǵ���o��}�����=:Ͼ�29?���b��`z���qӯ��FJ��+���c���zC� �DO��w���"�<s_��y���>����=���yK8~�t\��0e����Ƨ���=O#���	�t�%0��� �x��(�{:�k�
�v��?�߼�8�����ہ�o����F��#���:-�KtU�r�2y��Ң�e`*]D6WE�̬���Z���n��L�on��$�I�9]����\��>ވ����~��	�	��:��}�VJi�3�8�}�}#��>�_|�_,[��K�Pc�G�<xS�4�	�IC��
�\'����*fL;�ưa[7zbY�#Qh	��s�Ʒ�q��s��٪��J��w<�e�c�3��{(BS#��*��t"ֵ�t��e���p�هJ�B�n���X��ghnj��)���榳��ٳ�`k�C"����,߄�o/��KV����@���Kq��Sp�����]��o�7�A�L��0|>: ��ʐ�2�$�Ll&�kč��
S�m�� e�|��Sl\�	����c��$_�4�Y$=5�Lb��]ؼm�[Z1a�A�ӗ���;�d�
L�o.9�X�Q���ʭ]���|�U����6;�����1�s�MY���kW�t�!�9�4��6�M���G��Yj�W&�
L�0�:�T6I��ZZ''~��q���4g�0͓��	0P*�����Ibct�{W�"�*����q��.��~Dz%�I�5���a�D@e)'� ޽M�,N;�`�~�a>��B�?����.�nߍ\.'롹�	3��Q�F�^�B+��F,�J!,�y�v1�r����u����1l g�Tw��_{;���o`̘�8ꨣl��):�)*�c�F��v"��!:`�d�Qo� B�dR��Y�[2�[��B��ZxQ�	�ӆMx�����q��sp���̓�9����	L���k�ߘ\}Ź;�I�h�����=�=�6
h'M|�"po�Ko�E,u"gU,e���E;%N�hLe�r��45���/���T^�`J��S���s�Y�|�P�Ǜ��S�4v���՘�|�NL噫u��4F�U���?K�@mb�:/�^E����	�RF������﷚��������/�#^����Z'r��Y;�.C�n�=3$�sO=��~(���ۮa��"Xw)��?�K����w����ѕ(��
�L����)��@'M�S�k"4YK�4ž��e�����P��
Y�Y_�E�^Q��3�Y�P#�P�?��Q��bf-ԯ9qE�EY�#�����-�Co5�T�j��0�&���y�W�:����%���s�6� �0��o&|�I������e�r�g4�N#a�I�:5TPb�<[i��bh
Up��Sp�׏�Ǡ%�q!��[�J!57q�&�~>]�#O���VlG��$�8�?$ �����)0�ϭ�5s����Y��G��T1�&�\Ys��p��. �Yk�7��q&�s��"��F�]�-�*K5U@-WS?Y���F�m���m'�u��^���l_�n9<��Qc̐=��\��]-��4�J`���q�ŧbd�G�A��u�`p!Q^��w�}ړA�C�:)6T<=�bDI��T�[�Q�;l?|��s1c�Vuw6�g��P����������@8�n>zݷu��H^�֎T��J��S�;��c�޼�2h���z��n���0ճDe+0-��r���L�:>0��IV�9�>��4���� ӸPy�1�0���A��Py�#��9W�Pg*q1����	��������BA�j��d�6dLZ�(S�g��YW^O!�P�߿�\9� �ֹ��;~����j�]�
p�C���!O�0��o`��Ar����'����w>��K�a���x��[0|�Ȏ����#��	LM焏]���p-n���������9u� SL	f�p�kX��YP9�v��!�Ɖ3��3��ԉ#���x�ǞY�{�F�)7�@��+�9����8 ,{���	<@ӞW��k\�e�)�'>����va�i���7�@1�����=&��d�W���.��އp��܆�X�dRD�䌻%�ʇ��$��,��&4>/��!T����gX�u;R������b��arx�R��w/�6��*.ƸL��jtC�Q�ȕJ1�brN>f"~��0�Iu>RU��[ڱ��b\�����&Bettv��7&ο�HM͍��Be�ԗ���T+�l����4���ُ��<W}�LS�����V]�hE7��,���!V->445��1
��%��k�vT3qm~v�9����B��d�M_o����L��7�@*�'��j69�IP'l�\�{J���Ց�_�EGW7��2~����KO�OB�=2�����=��;�G��/��Z^ƨ��ΜK� ջS�k����Z �T7wN��m݉U+V#O"��K�6H�?�P0(���гY�2i��bhhj�1��}���҈y���0~�Q8���rs=�M� ӵ{���Z��{+����
�{ͅt*�D����D�eL{�Lj�^=��ʫ�y��F#2}s���6�9��oT*/5���D�,��򆃢w�y��g����׉� �sJPI3�6+`�����f�6�
 ��NL�&gm��9D@��dzLI��6���|��t�,���̓�"�\MΊȤ�����݁�H�>';��!����W�����Ew,	�׃��0�6	�:�MMh�L`Ś�ض3�\���0� r�?*E���    IDAT�Ĵ���٧��:-�0���O��܅=�X����w�8�0i�h�f�5�<��oC|�^4D�:t�LE�����
s��q��Ijo �h�`��A��}ﺵ���ÏJ�u�/�Aӧ��¢��?�<:K�~�����+/���M�&y�3���'?�CO����%wD&������P5wY�5�mU�ѐ�-���t�DV�ṇ�H�j���k��:��&Θ�H��Xf2f��bӠ��E�:�֐�Ni��1i�w�u�������W�'g��-p����N�dC>�L��ȥ,9��я�DXP�X�8F?�h���Q�Q��9�N�*�Nfb�Mlf�r6����<����f1	�y�2T.�n��ֵqm�&��A3��>Z�W|��]Y�f���"(Ȕ���'l�:�~���@o@i|*����J}u��v��,���RӺ��3k@kW31�k�Z�����2#�P��u��b�b�h���i�諫�M����*P�#�#;��0ͬ=�|v��!� u�U�9�)t`��身fM�/�
��Z��u�um�+�4$$��X2$�pg�#�*�؈�U��ȶ N>v�{�%CW2�M���s��a�2�agϿ�)���{ce�� >������ev��A����TZS�9"}���(D�D]��4t�I�m�J1h��V�Zw�d®YK϶�\u����g�B$���ߣS\�f�l�S=s��y�=��E��c�>q�y�e����C�N�5M��&^����E[��+Ξ�Kf�A4C-m��}8�rc�^��[�S����m��R�1�*�-z�*2�8�}���Cě�׏��_u!��O
�����G�]�{{=y�-��px�s�i�'�g��tn�;�/`;�q�C�q�)��
L=B�f�q���N?a1��(g
��.�@��N]#AT�[*��I&{0-��21�6���L�ƨ�?S��������%���K
|4�*C�e@�y�bɵ�5&����4r>Le�Q.�WJ*�)�}a������A�j��M������Ǟ_(�q0�0P�)�^>߁���'���Κ�;��1������(��}��X߳��7�?�9��;
��/���m	䙴Q(��������L4��	<Ė���O�/���}�&R��h��W���Q�:b?9cL=`<"�V<��G��c/c�ν"Ҏ6�q�7f��G(���=q,�`|��	F��N��<��*
Hٕ��HLݻ�g�*T�����³�S�U$�)lٴ�2�N�2�H��kF�ը�����ȑ�0e�)&��u��ȓ/��e���Ӊ���/��O8q������r�"���:�g�+��xiLdl��}3A؅\��n�v�d���1�Y7{y��@Wg�{:d�.Kƙ�%^�H8���F���r3$ЖIhX�|#�/\���4�a/N9~
�y��⤫�	��E`��{�ǪmY[����4�H$��ߋl2���6���ð&����y�D't��7K�����v�z}�'����R�P ��"���Ɋ��EW����vc��M�������}5.8�8x+E���y�����"�w��X��O�)i��8���:7c��m���aҾ���ȦTb}	�ض۷�@:�BOW��{�T/v�9��{��0`� L�<���'ԗݝi<���>|0�9m&��IUF��j�����/a{'�4
խ�!*�X�|A2ZI;v�U�{6�N�y�jS��T�5��h38n�}87�\�x�h[���V�)��Zt�D�ȩ%�n�%�2��u��@&�/"m�h���B��B���h.j7�G��q��:�F=D��L4��R�5��	���Śd���ȥ{��)���'L���:�b�$���W౗���]�V�8����s0vxT�&��Y��=��$�^ ���FeP���Y����ְ6�jS�E�{ڻ��;��w�a��'r���ޭ�E{2d�0���h�hT��'|�cZ��w�A�$�U�CukV����܇��G�o}#Fs��d����_�'�~��&ǵW^�1C�z��O-��O��<��T�`F��P𭩖R�5h�SA-�0a����l���B*î-'����{Ր9�� ��b�Q3o�U�c�o�J,�)�̡��$��N$;���������X0���R�'���z�&�8SKk'�N*�k�}X��4����T>��"��Y_�ΑԒM�e�I��G���<%Ⱦ�2��Y6;c�%:1�Ճ�f����¨�@��#sqE�h���#NI����U��ڢO�����ۀ�+ 7']F�F~eu�ܣ��o��R1m���z`Z?1���(-M?l}�oj������|� F��l�Ԩ�4=���}6*�h��a
6�+%�+��ez��c����	]��2ٵ2����|s�{�>-��Oi��Z��S0�Si�����jZ�F�i�(�7m��m�*�����*�Y�|����Ǹ
qx�)L�0�_xfN���{6���h{ʚްF���?oǃ�/���=(������aT�f)f�ְϻ�8��V+��ka~�֊m���-xT�P�:��X�f�m�Ѣ%"N�ϴ1l����}��j{��&�~Y=�}����hX�k�l�65�s�6.�b�#�c(%�y�%��F>! �ٛ���K�:F��TS�zJF����r�kB�E�U�I�m_F��g(UK"�J�z�\F%��+����k/?FE%�<��12&�Z�{��:�eچ��(9Ԝ��YY�{T�d�%F���P�g���Q�?D����O�A����$�x ��g�U���91��#�����P_B^��p3���sR�S��C���T���f�	���r��67��[e�ǘ/�f	��`ͯH^�v�9�b131
;!-�T�@��+{��}�$��+ZrL��$B�|��p���f4���3�˹��J5o��m��ǟ_(��3�1��2<A�=i��ђm��`�_�9�pӯ~�ɚ2�R������P��	�W�{������]T�"�s�<����h0Q|�}�>�?�7�&�ձ���2�?|�<kfL� �/]�7�� ��nB<އ���7/;'wB�0Vm��?^z�.߃l5
���/����� V.���
����؎�ͫ��t�o���9\ctL)P-��RD6K@GM������B�D"��j�l��S�m�����:0y� �q�/��4p󽋰����#��R�j�NL���ƴT�#^��.�z�$��rbʑ��=J�*r9�����k�͈��L"��S/�S��8��Rh��9c,.��k0 ࣕ	���+ذ����QҡQ`D����-��m��6~t�8m��������ڵ�:�Ie��ك��N$�I�y< �GE3]]CA��yI�v�N>�x��7��Ͼ� ���"v��~�9�?հn� ӷoǝ.@w܋\�4� ��L��n�I���qȔ����1~L>!�s�|�-���Cow/�zb(d�'Y�..͟[��Ҁ��� U5vu����0|��}ڱАK&�^i��^���,6�3Y>�7����Ԝm�4����j�Gޥ�W�	6cI�e�2sL�L]?1U:7��8qrz�J$ilB���HEё����f6(>M��-�*YL}����ƔT^ۼd�QNY��E�Pq�S0�LA�N��Ip��,D8�/�ޡ�����Fؓ�Esf�ҳ�HJ�[�� ���N���s�w�I�x����',�an¤��n��E�\�	xdoa��P̢ZJ0=��#p�UgH���Hu�A���O7�b),[�zz�0s��2����5�[ʡ�}72�� ��0j\F�Ħ$:@�'�.P�6�Qf\N�?�K�,ŉ_;L�� �����T��%|��q�>���`���zrbړQ`���� [iB�߄*"�j�/�Aԣ`��\�Q#c�>��Q(V��������\��ƘEM@L��q�6ۘ��9����^ev;��YW�:�޺`t��fZj�ȹ����q���a:qV�i~��s��ze:��n�i/���jtPuT^;!�i������M��X��8ѳ�L��83�1��R�\��qfJ�c���"�� Ӌi���S���'O��41
SI�:y�eA�,�%ݺ'��o-ŢW`o_Ep�F���&��(�i�M����h���s�Y��.�b�~����=��C�� �|���kfZ�Mu�G�]��wic�������8���u���w��j��Y|���6��4�����3KI�0[@�����QV�V��ʳ��A�^V?i׾���i��Nt`��l׏�[�aHj�S?�46�XE��+Ҕ���R>�R6�r>�A�^�|�T�9i&���Ҏٜ.R���-21ֲk�V���o�����(�w�Qr�$����!��~��o��a�p���6���Y�kv}�/8q��T�Ag�f�����2Fj�jd:eWa���*}�i*9�x��+3��1�Ss��v7�`�D���ƊLP���ʣ���x-8��f^U����n5ۃFO�<�k�����ɩ9��R��Kz������m�p�%���|ƙcȼ����<�M ��J1D=Y�<x.:�k8������������/��ɒm��5�LG�cuZ��'����,�����+�׽��WA%c?JnF]�e`L���e ����T�+O0�đŗG���/ڀj((���f�����[s��G�)'�J�%0�"��4��WY�QW<DL�Tcdc7YOy"a����	�i)W�m*
�Bt�&�ϳ|k��$�PcJ��]|2�5���1� ��e<��[L9`,~|�%�1Q͏�`�g[���ƪ/��e矄�����ÿ������6��������*^s)���EK��H���G�7?�TMo�k��u	�r�kذ���8��^�}L?�8�8�:|2��������+����<�ӦN� �x�@W���j<��blmO#nV�B����Nj���;оy������p�Y�;S�˞b� L'����>ߣiڙ�C�9�2���?�g_|{��}�?�7�D*����k~�B,�p�Py�U|���腇QE|��[*�T�`�g�0?��%��lj_�g|��&��&�r"E��dh��x?�����+�cǮ�8x��=�5����ū����W������Q(�h 8����¶���ލ}�����a�xZ�B�e����/��Ƀm���Ui���Z��)�h����5�����a�D�>��?����p�����jL{S~*~�#���� �C�l
�x��q�����o�}G��@�v��n1�9C��q��ᣵ�T,��BͣY/�-s����/��Q#��3g�X]������w�`�v�x����
���ȩf�tY;��"u�u���UX+U0�>@�LW^f��#�t�X��`󆮰���RqdR)�H�u��:���o6������O���I�ͪ+o��C��	�A-b~T�����R�+��x�:W��;�j6?��f�Ia
!�쒊Y�T�JT;��t
���7ď?��;8fz��A���8���_b��Ո�s��8�i�{��R�m3���?��-�70�_����J�>T�8���p��:�uf,v�c6T[h����ݎM�7a��1>|X�9�ʜ�"��^�vw��e ����F���V(�(�}�(��^�y���b9|��'�`8�����л	L������������\:��A�{��1}��%��s�!]iD���& /�,�NX�&��\Ӷ��1|� �&R��� �a6��:8�1��p��,�)��)���	�eH#�\Wݧ���AoZ�=:�4kf���E����;�	����f�<3Rw�y��Bh��ŴXGa�C�r'�z�1,��:��I�uo��Y��*P�?��W<�L�m�s���C���9�rq��I�t�$�w�1�6q�Dʉ'����}8��>�7���Z���j��ЎYR����-�h�&M3��l,��ժ�3;ŢS�������n<�����R_-�r�	Q��1�ƅV"���8��z
���5jR��`�',]�L�~���NAk\�����p�g�4k�-a@�:R�݊<����G*�1y�	�i�f�GFOZ[�
���Pg�e)�֤̮aEG�ss��X��)���~�`H� e��3��:�&Ľw���8뤣����1zH�q�V�i@�	dDh�����3�c��<��(y��ƘAP���I���ձ�,H�ur�<7��-��i����B�cW��L썩����οP���i��'-Mk���n��i�|2+o��߻��F�e�X���u�l�2\rm�hL���٠N���C9ݍ�P��4SFCFOo�����[�iGU_3\|�M}����"Jr7���(�He��Mu�WM#�+c�A�>e"F�ƆF�}�l���wWb�^�<����-d���kbe&Îӹ�3lȳ�~�{�mވ�/��/4\ʲ�{緩K��;��-��O`Zȣ�͋�Pȃ��"�F�pE�"���D�/u�:�V���)�i&&�&���ԋ '�̍�)���Y3��q3���R����I&5�4RWߐE��F"�x��Hp�&M�DjJE�ԘFʽ��"��`?�_�>����^�c�/|�����Us`�؉�>ڈ��� ֬Z����?���L��U�N�Ǯ�H���&G�������ϐ���� �+������|��JZ`���n�|��ظ��\�t#��������هaD�7T����I-3k6�d���8��e���"|��6�\��表SSd�*�_
���ۻ�7��;Ӊ���E0c�´���}�Y�U�+BĆ� ��փ��=��z�<�īx���`o{;�M�����>e��Å�,p�o���둯�QB@�i @��=bܤ�j~ĉi��N�9���be���J����,��.�bH(�܋d#R*$�9��+o.��у&Dm���a��+��װ����!c���	���&���c�Z�c�����}N:j�S�\��l:�	�&����{.w�����uZ.����n|�����X�|���w�c�iG��*���	���ۅ�ۛ�#W��C粠W��si$�ۑ��*����ƍ
���B(������>��4�,4����ޝ��Ͼ�Ç��3�Z3x.#|�v ?��	l�SD�9�l��1F�/k�Z*���=�l�n�$Ŕ�LTxg9�(�� '��0�n:�音�p
h=� ��qy�����\,nt�ֈ���:�rbZ��s:-�G�_0��S��0���'e�P'뀿X��|4W`Z��`����;SF��)RDs2`�iRxgR�ܾ�O�?��8p�W�#��r�7>m�����-�H��]���P|�0����J�r�}yi�F���(�ZA! M���,*�8P�Ĺg��>SL�t��n���6, ::��Hf��� +�˾��d�������}qJ.46��Q1���Hhmk��Am�I��  _SXc��lݎR�����p���ڔ�>l�u
0}˖}��3�÷.>�2K�Lzz)���{HUubJڰLL�XA�.��ǇY�!A��%D��^1�5��`�^����N`�r
�B�RX�e6c��z��m�֦Jْ���[k��"�t"d�y;!���)��Ҕ��\á�ƽ6�jٺbS�_�k$uŴ�qڶ�R1k�T�^'��&�Т�R��כC2o��K3�B��l/��p�iG��3f``$f�Bq�k1I3�$�b�<?�=,[�[�^3�H)�/1��6��z��,{��ɚ�[��z���ɏt@�i��θr�� ��	�W��\79G��Pꬣ5�YW�ZdN"�0rq*椃rOb_�B^�Ǖc4��B��9/�Dy�gi@�Rd�B���!��r��T�N"kӵ����6����>b�#���5���d�n&�����.���I蘉	��BXe8�WJ�6��K��D�8�H?J#�<*�,\�<*�>��8l�X0�Y    IDAT|g�l�<t��&��o�&t�w�1���I�����Ξ�� �>�;ӓ�g9��f��hɵ�B��:￶���]��r�^����Yd���I2?�z4��S�ZݷY�fo����T�1��W[h�͞!���~u�ݽ����1b��v柡��%S�!m�/X����J.&�숯��� ʅ"�,�
�0��6��Q�C��F#��
��|Ɗ�)�@�`H��B)�|>�l��\A�!�͑��~�=A�>$U�4�	"�|P���4���bA����?����y�>+�[����A�N���H1�����\�
�e��H�Lv�Ȅ���b�B�<M���sڰw�db�J0�A�g`*��Fc A@���{*/�)�i>G��O�i�1�
���6�Tښb#�|�b	�LV�)_?��1�
�i�	mN�w�'Ĭ~���sbZ*�[L"Z��w�?ߢ�/��L{����}O���<���t.fL,
��;�ǟ�r?6�[�����{o�	�a<�����i7������kx[IAd��x
＿
�5!^>O��>����&�0��o}���5l��#D.Ǹ1�$���G=*��h7|�\R�f�)u{Y�Wb��
���'��]�����1?"Ь2Ǵ����ؽy%��Eg!� zb�6vS��?}C:�3TK+�LP�B��B{_	�>��x�e�޵0���1c�8�.�h�n�}��h=2�ʮ B�����4���ʹit®c��B.��O���}�"���2F�jL$xh�Js e�\2.l��N�"T-���q;;X��FlX���,�7'����{�wy����|����YEt�y�����y���F��(��Ec��ל'S�����DRP_��M'U�e�����'���q�3���a�;��*�������HH	��PQ:* ����XFGGg�u;("���%҂�Ф�P �ׯ���9����{���D���x���r�=��~��k�C(z��wF���^\�*&M��{��2�=�8��3W{v3~��G1�gE4���d�(��Ydw!;�G:߿�*̛�b&���k-h�$T���
Ie�UF����[w��+���,�@o� �����GF���ad�)�U�4"�6L4[�g�2�f7`j�5�� ��.�.�:	�I�C~]�P
#(��He�ŕ��E�b�dA��}�2�Pui~T`�_�1�ا����MMW�
�X��R�˃���q�)�>ғ����ͬO��c�pC8�U�/u����]������eX8]�	w�x�ͽk�[D�ʅ��(2q�� ?��j��&L�Q�>�?��A��.�B���ɺ ������? ����`,�sK�]-_�G%����|�7�!�f?1G��zC6�z����Ob�H���O��	��4̟���<�.Z �Y�V���v��1U�z �;�P$cp^���5�-[A��\����o����ŧ/�fO��X(2��c��;V�w>�b���¸����[��7M���}��k��-[����PO�(�E$���e�s@�!�<��$-��:�	�T��4��ug�c�56Q�Wtq�=w�9$q��+{�:���\Џ��&(��0`n	��PAbksw3�q=�N�`4��r��-)���d�d�ZF�2�L��C���K/8	G.������CarT�!eI93z�.�w���5 A���}qDc�E�]uB�~pc�p����S��ZRh@�"Ph�M�N�]+0�~Ka���o0�)+�t�����cg��<�G�o�>˩k������[Rg�E���v��K���T
��z\�Z�67b�!�.65ע�ae2,��V@$;�{I���,��*@Ti2�c|��h#=�f�E�&��z�V�lF�/�)ڀ��I��;C3���b�sg�6~>>���h�C~���0z�\x����0oF\LphB����N��%{�v�����<�jJ�D=̹ʴC����a����X���\�ȝ���n��;�+���\�%���Vu���9JQ6�M$���Ri�@
�L]d1��nϽ��{ �[�Հ3QwU���!��\�[�\P��x�ʙ�V��4��
���Q�zrvgQzo�� �B2ݭũP�z�x%��%��7���*Υ�[1�F��Ea��zѰ�X�*��a�"%�40�B<ݍD�]�)8��`�����Zȑb��Wwf8����rŜ�(���M�1�	0)/s)�kA�=�("f~�!T���Ǵ��W��(�e��Jyi��h�sx�Q�L)�yUx��0�t�u6��b��ZClv4g�R����Qab_Ig��H�T�qMR��Tn�⛽�rm|��z)D��_��G,Ӗ�)=��%���Ww���=)���\��?	�.�"�T�<��&����7��e��7��;iS�*�4���&�y����� �����V��j#8j���Z��x$��O;����"�`Z�|�?���ذ}�L}��kr�]|:N:z���&P����;�xp�/�d=`�X�
�o�kX���d�N32b�D��,��������4\�o���;�0iJ��h���a�k�L%>��V�̍Ƃ)�K�d�*:4��W��u�ߌU/�.��e-���/8�%�|��]s��x���(!�*�H�Rj�T��jcL��V`��ʙ��e�B�	���O����H$O�؇�ʲ����s��ҫ�V�Ĉ��"���.���p������(C[[�D��a�o� �]y�}�%8��Ɣ�'Ë9JB�jh��;�T_�����q�?T��>�_��l޺�z2��5�����S�
�th��q�o��l9��O�"ɘ�ci�N`���h�Fs�|��{Wc0�"Lj)��>�6h���F[�u�o�����mø���d&�٧k=�4�����xS^-�D�Mf�R����@\���4m�;E�#F4z����8���/V�E��X-�!aLke�a�K��vOL	6�&�
F�4��UV���SV�&���Dj���R��S.O�-2�$0�r\��"^�C�`�8pj��<���!w&�|T�c�m©G-����I̦
�� ��+�ǯ�D�0Q@!�C2AG&�Es�����fw��=�	��y�����l���Q�� @����ӥ�����4�){�O8���G�����|itl̀Ж��Q���}CH��r��:�|��ڰ��E�o�>ℝL�11Q��m}����/b��|�gb�A�����1{gY�ڴ���o��6n�ǎ?�u"fL"^���4���֗p��Ϡ�.���0%0u	�&{�PA�E�Z*�\�
�ȫ�D]��J�B`����1�v��T����q"�3豷k�B��}-#[,���2p�<�7�������+�8`*��%;�|C������%�D6�qn��޸ww.�A�.0�1�KKđ^V>=��Z�(=j�+�y����	������sc�ܐ�gC���x0.��c͆,�{��x�ghD�K+;�SV�=��[M&X�HʬE� �W&B=Zw�-g`��9Vʱ��)zG[���
}� x���{k@ X;��`.�\��9XC��N:��:G��!��Z��xo���Jq]��5���׉�%��A�ǐ�C�R�C��D%o!���9���],F*Ό��*;��FM�!�Y��}\���/�Hq�lr��e��)���]:�{ֶh��Ln�Y�b�HP��a�����B&R�X��N;�,���˻xep��&�!`� p�#������bLZ�wJ�7a�e�9���������7�I�	F�so]֧knpjLq�Y0R�����RN��8kY:hCqlk�����,#C�V�U-칎hER��m��ɽ��>�Z���h�H)�,��Q)�P-e���
�x�,���vw��{::��<�0:^�om��7�b��@=������{u�S�K� Od���HF˘3�K��ӻ;�b����o�֝ މp"-#	cI��G�A�{R�87�Λ--*���P�Ń&1��8s"S��!�)~�������P'&�=�i��U�sA�hE	����yU��� S1?
�Dʫ�4"&�dL��A`J*��g�3�jܤ��Z�q1��co��r�AY{L+~Q�m�'""�ckZ�>{g�fv�2c����#�e������O��ӱ�{��-�8h!���b��d	Ɣ.>��F\��?b��o`���p˯���;$�Q�M7DK����G�A�ɶ�� P��K����W��w��5ٌF�O��y?
���y���Ԫ~��懰���Z��|n!?������gcތ.,=`Z2O�E��K��d��ӂ<��j<���vl�6��D"�!�q��f�@�(x0��pl`vm|�� ~�����:B*�<r�{�n�F����OE`�{����r�2F�9J�=�/c`p��l�sϿ�g�}�BI �����O�|����X#c������3��آ�26�QC�+�L/�JyM�S���m[�l��o �-��l$VU<Oz8���dQ�>k�̝7O�N�)T|<��<���90��6�v����׾�N�ϙ���0�~}߽�V���,��N��X�t�D��8vl������p�G��͹��$��(۷�^����]�+��'庹Bcy����)�)��X�`ݻ[q�}+��s/���bʴv��5W�O�9�L h��Г�?<��R%��D&�H"*�hBI���}��.>p�����sf��y�t��1�Α�B�EΞ��W���p��K6V V��6V<��o.9�daLU.��t� �k���C|�R�Ntww!����ƞ�|.�J��y�U�"�ǙR��'!��Q{�8�U)�)���j��A+���U�gab�b^]y����Wf`�D����p኏PQ�6�Ҕ'��D=]h�b2.�����e�PFD{oxv��1ά�����Bؐ���EnpN9j|��`n��/f����W��C���}C���@4����8��}p���a�����>�7��8��I,�K��s��?�Pu �R�{�i�q�K%�
��Y���29al���;��ۛ���w��yJ�3U��zux^�D�tFM�xp0����:3i�	��Uq�淲�,��GP��2S���O^r.�)�[�\��K��ol�-�-G������sO��N��l\L���U���+Qu�iG�U����1U�eL�-(��ƾДo)9jI�J=�,��jw��{��vX��d]Bv�%�M`��c4�E"�rn�:�U�nu����a'�T�(u�U�}�Zj�II��U�{$�R@i�7r����[�,}�Ĺ�[%�dե�����O��S����B�tǊ8��C�OƬiV��Xb�����K�}�ҚQ���n�0
^~� ��q)#�L���!%�fO�1��.��$0g��T[q3�l2R��T �k�����l�:�V ^b"��)�'d!�����,�f�����)
�P�=�l Q�F{8ŉc=���g�dY\mH�-#p���
#�0{#��ż��<�!�(E�)�����\e���1��j�^��� �I��V��eԓ��p�j�ɫ��w�Y�n�~�R�+*٪�Z�ͺ�D2�&0����Ĺ7��1\tƇq��G	1�v.�qT9��a�,�d���y���1����vY��/"���{˂jP(rs��Jj�r�4�bcԜ���7o�s��C�L�fa�ͭi��:�E�̍c5Cæ�R�����r�{6�0���*�r �֝��k?������}����&$�����r�����r���e|�gMAw��@�Y� �vP]������ݨF�e�D<�f#Kꈧ���/��ja��t��ӏ��:Hf���e�闶෷�Į�**`A�)6���+��r��>&��h�XM���݀��\�Y["����E5B�(4��~f�}�$��T�>��WYzL��F��)�A��'<S;�5Șf8�!����IV�D�a�G�R^�c�g�B�DZ�k���^UM�MdL�Yq���kϠ�����z�X!�z�����-Sʀ���#�e�1���'�sg.ä��1m�#4?�aŭ�>.	����W���O��Ͻ�	?��X��L�����*N?�0��x/:�U����r�ͤ��g�P7��/X��k(U�xP0�����3���|�<��d��zi ���Q��dh`'��;�����8��\r�Gqŧ.���v�z���������>��j�ba�s�H�sA���Pce@a��a�ý[�K�B/n��|򼣵5���ո���n�v�]]X8!&O��d���5a&v��C��=~M�Jϫ�\����b�!�4�h�9���?�� I0�����ɗ��T'c�@<��PV2��/�*jU�1����)�7�xf�3���0�_���v��d�C�ZUn �x*��7�ոg�$�|o�P.cxl�rE�==����������͇��;�}e߹�OX���D�L�	<�TJS:ݎ�mC�4�)�*�u�8��K�10ǃ�8�o�V�|hD��g޼9X�d��@|�ߌ�׭��DNd<C��q(���q���Y{����w�����ҕ7�bx��u��+���DB�joG��!��(�<��v`x�:s�<\�ïcެ��F��7ּ��+���Ξ��~(�̞.��1Q��l���l:��X��s/����y�����o?\�ͯ��+)���.����;�s$�H��.ώ}(��R\�[��5�`=`��tW�&�늓f8,=���ĕ׆.�I�J.�8M؄�8���i����J�+/g{�TX]y`ʏS���<�{V��� &�َD��q��1UF��h	��C�\Ce<�%�A�%KL4,�q	�D�LH%�AY���������ڧ���j�d�L�����<:^3��#� ��-��,�������o�N����J�{q�j?�;����?&���d���h�� �\��8Ac�����h��R��B����a�����8�&��GV%!�l��害�Jf
�GBȤ��𽒸��rèW�Fh�T��������n-���ϖ�k(���6c���V���E�㲋?�)]lPfy���m/ʸ2��X���Z�Yr��l.�,Rٕ�6)^ݘy>����<��Yr$&X�	nJ���xk ��J2I�9gXt끭L^(��ğ�9��~>�`��u�3Ry����HM�/,�K��<5��@�H��sBu2Uw?�e	WKy�\'�0����}|;����=����,v������L�X�ٰ��{~{}v�z@���<�p��19��`� �ڜ��d�����e�h�9H=$�r���.E�	��/՟S����	(5Ŝ��^TB5)��Iӯ������AdD+�4|��Ue|\2���і�s�-��֊D*�X,�x� R����]
X~���g��I�c,`��Yo�P�P�jȗ<K�\j�Fԁ�瘚I�̑���Չ��Ɉ%R��"c�i���vFz��]+�L'c����p@Әl-����jiSG4��)����F�4��d_��P~��.�>�R�Z��0�By�t�����Ӱ�N�٨
2:n�R�Ap:�Ͻ6�_��^��8�j���I@�^:v@YA�Ⱥ�R��Mkh(}�N��$l�;�KP�o1��_2S���Z��� 5?zo`*��E�v�k�be��]��6��ɎT�9�S�=�u5�r���PDm�2*�a�
�N'~�o_��}���҇���+�$��{�]�q���0��[|B�����l2��T~�r#@e>b��ٓ�tQZu��<��m�������[�SHut#՞[��_*ʁ=d��0�sI�bJk�0���1�s��A����v�c�g�33�
�)A!�8a�%�NE��N�"mi��BO�8�XT���)�t,��F��J.���+�(��m0��,��7��K�y%0eN_(�\,�ޏ�҈dRB�S�ڥ&��c>AA�ΊH��x5��7�+�;W�u�Hy�E��B�F�ҕ�z*�/    IDAT��V�9������J�)ߗ������o��k�!�(�������	��I;�kY3�%7����%h��([*a�_����p�o��������&�`�q�u,�q���I��L�x����Q􏲢F_�6њǐǌ�N��R\p��8l�a�4�V`��H΀ޱ*�|�E���*�JL��+���DU(�xН��u;6bp�:��1����?L*tZ��T����+�_C� �FGt��tJ�
)O��\|��HQ��&�V�ˤ��;o6N:�C�<)#��z O)�Cxz�V�I��I�X� ��0{^�lFW�J�B/�8~�˗��J�esQ���m�x������8��%NLV(��-m�}J���H";�t�r	�}��Z�m�3gN>�CXv�u,�����^������*#�>M�8Zn�3$bQ��G��G�4�������q�i��\<K�F�X���x��WQ�T�yUtO��R2����#����\�^�dm�6h9C�)�/��+�K/=��?b���ց叽��nY����_K���t���R.`x����Ǳ���O�Ϙ33���]������[���-[���<{Ϙ��Tc��+ȯ��N.WV�Vk`��x���a�F��ęg��o~�*�t���x���7��vUPE��S�L�YV�s�,JE2u�pX�@R��~&�D��B�ŴgkkC�=&�*��<,�L�Ji����(ʥ2�]�tw0��\T���D`J#�H�\y�ԋ�ˬ"2��	0�O�B8�T)���jJy�I`J�J���/2k1d0�$zҪّT���v��P^S)�<я9S��¥���EO��&�hE��EC��F�������;�a+�=�E�"�+���f�p>{L�8E��%>5�Ex+뢊b���*oG������|��G���xl��X��u�!�����ec룉о!$�qT�;X/"-c�y=��ޘ={*:2q��Q��3��Tk�ȕ00<���q9��>x����EHs�3�������??�2z���H�w �|B{g`s�ܱE@�l�V���9�B](�,iMĜy{����V9tp&�� N����D�����Q]4���`����	L+�����B�%�p2�fk%ڽ�;˝�L�"����㯁V���uB g}��H
�G��K���(y��R�̨)qF���1�3=��>{&>��2:N�A�2A"�#�q~d?n��q���Y/�x�d��qY�|�X�Θj|CO{t��'��6�k4���BE)(
�c뱔�H�3���
'�k���pWKo+_��-q�Ws�#��c*����r�O���D&���:���H"ڨbrW��ľ�������ن��6$��j�(8QX���)�V�lI�ma�	�;���H�UX�P�T����X��Z���;��h�|�r�
' � lf��La�%��uv!F���K�8�h�>�@�����&9SAg:GW�r�E#YK���;k,'9w U"u�����ع�:� 	2�*�gg��E��4��8p���O��;�,����\�r*�^|s���	�z�~�K��G2sc�D�h�Y�T�>k�͔.$	�l�+���~搎1v��ڞys<�2�f^i���-)���kw)�K�[��q�VG0�����	n�ˊ��n"��MӨd�Q̲���5�P�g���B�i�W?{6�Y:3kt*?\�fa�������p���1^n��b�$"����c��
�HEJ��q��Ϝ�E3"�c�[DP�s��_>��x�Z
ṁ�u�8ZK/��N'E�y0�`���y>X���[���2�ok��,��Q eט���������Ȋ�+0�a<L�p���B`��G$o'0��E��H`*Rܶ��1���2W�X(��:�l��4X��l����@q=��`�h �����j���T�!Q+0�����3���;�����=)��Ϟ�C��&7�X��v�'��	��mF�/b��{�߾q�8l��t}#>Pm��rEk�l��*>e��=����}���P$�Fu���a\r�	����+��z����ڛW�w�ij}�P-�`FOW\�1\p�	�>9�|
�dE`B H�?VUv�w>�2�{�M��T#�Ty��Y��k�۾#��l���뿋��Dzm��S����EGV9i.��)�Z�,L���>�L�΍��I�Q�jM�O)�$c�������(�lg%V{L�߫F��A`*r�J��ӯ]y6�jәF��Ɣb�Ǎ�}Nb #ɍIk�`o�7�h���!Y��w:�D<�}���*y�g_Q)������FIYXJ�'F�0>ԇZqS�������t�7&�\k�G[�Ÿ�@��%�����(C����X$�8���0I�b:��&�T�0&��_Ș��8J~;*����D�H��U`��.>|���?���3���=[���U��7�R�^�aά��g�|1%"�+}f��T����7As{{
��G��=�!K�.F*�DJ{��PE��?}����H!����M�p�\^�j��&D��E2�s��:Jy|�hKKЭQZ¿s.�w��K�A�*�GEL;&	0mp&�����!�F'Q�u(��l|��Y�{LcҌ���#�!��tԓB���]���:*�9y-�ϫ{�_�s�k�~t�5aOw���D'��a��6|���p�ôMr\>����Rl0J]i�����C����ϮA�K"Ls�d�r~�C��E�6�O?
_��	?tм�Z[��� zfZ�jMBXj��>��_���|?���՝��:13T�-~�d�)������btw�	�0wfBh۷���I�E
%s�5Nɴ�z�yM��v&|�F2�w���?�A,�~���Ce���p���ޫͽ�:3�"ޣ�,�f�80�u�}a�_"Qz�����z�{.1�ח�`��;�Di`fB�9͡RMjT��4��?�"�7��<j��&����VF���h.���u�z�S
��ӎ����1��S��5��Ӑ#����^n@����i8���hg�al�`j����V��^܅[�\�����qfd8�H�Mz��9�Ѳ3' ���A��C[�Pp��p#��ۿz�X�ԗq����*~
>��V&���B���j}a182�\̋9I�R�_��"b�z:Ә7w/,^2����3z0}j�8�v�%0yR���ʳ�ej?�+j4�����l4'6�Ɓ��ߵh��E�%�#�cx$���,F��(ɟw���-}غ��c9T�4"I ��P,! 5�с}	R4���XZJX45���07p�+5��H�[��J������9`"kIћ�L����u�z�\矮a*�B�z%�8�0��]|��g✏������� k�`�͑^on����zO��Y��Z�L2c��f頻4T��� W�=��)�Z�����f!Ȝz��o�ݻME�.{-�Ӵ��F�4�d���J@�.MP�X�fhr���	�J��y��P���դw����3g���Q0�W^p<N9j.�(�����up�n�Ly��N�c��V�ob�C(ގp2���Q(�11<�ji�~�0\�����������1�7<�叽�J=���HdRb�O����R i��W�[���8�:a��#SU0FRI��P�Ts'�~sj,L��P��ע�_�3Q��j�0m� �
�lc�8��cg�J$������@�-)=�>1�M��s��x���8�t�'�JF�&�	 �Z��)Aag,ׄ]P�(��162.�Z`��q�ʘ�q1�ɘV�Ն�`�
�������r�G/�_��y8t�TY��Z/����p6��	??�t��E瞈/^q�O�+kj���:8]5���ii�W{e��׷�nّG�������-!Tǥ�+0%��/:�=�]���+�7Z�ގ��L��㧾W~�dLg����Pe�?Z��k�cæ�8�C�}�+�����:|�w��b[M��6�[ �Bʘ�lGnx��q����C�Mk��qÑE&�*�Mɂa�z�a��w�g��D�Ur���?|����Қ~Tji4�iD:#P]�LJU����UP�؎�O>_���F�(c!Ě��{�"�y��ۗ��C���� ��r/�	�Ǽ��韰y�C�{��UN�����"?>���Eg���ҹ����M��*��o�Qz(��9�S�������y����4���F1��ɣk�?=	�э|��D2#M�d�z�j�Ў���߀��?��Ƭ�qS�%�"�*��.3�87Mg��\�et�0��d߃��p���1� �ك�~q�R1�����^݉�G4نt:#`�F1+|�	���K*�u"R&$.�b2�GXIk���fVˤ��	�܋�{E�PD{�dd&MB=SC ���d�r/��iH�CīTY��l�"�+���ݨs�Y(,�}�Jr�s�h�C)oH�ŔF��R�"�ᒘ�X��	��[A��\Ag��{Di��WʡZǔ�(�[�7f�5]m)$�I�n�7�'�m��:rE���l����ME�dP��hK�Q�)g��rhgqΩ��˟9Ia}�H)�k	��:��jlR�������ߋ'�]�z(��H��{f���n�IA�y�QĲ%3p����}-&L�f��0�� {=�*���) U���:~�S(T;e�(��gt�֥��
*}�J���y���\`tT6~�f8k�<E�V�[��Ig���z�ZXt;y����j�i
��2�A?�mo�)(>j?�|�"�{ʮ��N��Yj�j+�i)f�B�|�xu%qҤY�1O��B�o���gG��߀�{��+��'��-�hR��ly	x��M���簹7�j8�r="1(�ٵ1J��#�F���#��
�-���;6� ���A��H��ĵdS�**L9��3V�� �h1���(��,^hT��hJw
�;��3����s1cF7�x_"L̓��\3�m=[Zמ��`�mP�v�۝Y{ U��-1 �
.g����k�k��B�"06VA���X�O��U��f3�FٛN䐖�@$Վ(�S�#�J � H%0eш��:�.`�$�=���T�"������ց��zЫk|{�=eo`�Q����F���W�W��W�����"]v�ɘ%>6�@d�U)���-;k7W���ǣϾ�b5�h�[�o��Cf�;��~(�eH]o���>�k�ڲ�I��?�{S���RS�XQ�]{�2S*I��J`�f� �k�*�L͚�:'S��j?�yTC�aV���ݕf���+��M���D'p�%�༓�����D��WӔ��=h�W�G�j��~r�}x�ɵ�#��2��.��;60�J~ �������O�yS��"2f�,�9��W+��)d�� ��5�5L���r]�T��R�Х��5ҋ��֩�?���`�9��vԘ�lҀ�Pu�w��jɘ���Z6)���@%�J".�O:*Fז�^5`�ȗP�@��G�cF���L�zR��4����-�x(,R^���1%0e��v���DTF��y\G(�-XR�heٙ�S,�j�R��U��TGq����ʳ��x���� �ݭ68�=����ǟ�?)���/�UL��M.5�xy� ~z��x뭭h�y�����s?~<�����ө�E28N��������bI��'E�U�[�Y����zK���ك��`�S�6��.9W�L1?��'�֋���F8��Jy�<_���p�< �xÃ��h��'_�cϯ�;���G�{?>��8�g������X�v?��n0?fa⩖�zJpQ*kZC%?��]����׿�N��^�l��d:���%l5�����\�jOS�1e#���ן܅76�«e`�^0�3j�P�Yt����ѭ8�E������NS��$YΤi���V����Gb3Qv��s�D},F��S.����nG.�x�d1n��b"�:F��G��n�\u���������rWq�&1��q��{�����"��1���U�4�i >�.~ۓ(x ��� s� �݌��v�|�|��Wa[U�oL׎0){$�j���\�ns���n���500H�c��_�V��^=%s��ɤT�ݼOwɾ}`*.t&��#��ʍ��kR^JTL%��T�E� FǼrűQ��Et�LE��[����Q;;ƚR*}UԲ���@�l(���S�PO��gB�T���P3`�@`Z�`�Cʥ8Qal���
<Z����u3e`�$B�T@�ZF�^F$��`�8.=ddT�Ƶ@F��a&otL#� ��j����8,FT*%T؇���yҡ���'��-3 v[���=��&B�����=�GW��P��ݳ���\�U�e$QqM�wn����ȃ��0.x]�{͏�R���F㟹�<��{����~;ʒ��2�������6%�f��	�eJ��P#�t�Z���P�_���RT��������.�٦)E�뤬LǀJ�@�~��"��5	�T0U6��&c�c�»}g���uЪe�F3z�y�w���5�M��a����~M�Q�l{����9��:އ�u�+�;'5��K�k1mSY7�2���Q���<��y	�j��$�T;�rp������K�p����Z��w+�������9�I���R��)�zġ_a�$r*e����r9;�0�h�G&��i�p���8��p��0{F;��.���H,;#u��}Yb'v`¶�fqOT��^�7&8�ZZ.����V�
Q�XTw?(F.J�F��6^_�+�ߊ��q��+�E��&q:ЧM������)�%�Ȋ�����Z�h�d��ZL��b��TUE��o��m4��f:`gɐ�;�o^�M�4^WK���&p����<.�� �}*��uL�ds?p�=\�/#_K"�jGW�e�E2�J��|k��3��Oo�1���8���ֲ�[㺈m�X���q���}�M)���[�n;�RM����bĥ��2��řJ&��2��<W��+n-,�����X���H�q�ǖ዗~ �1H��{�-� |����
1g#�1�߲��O���ע����1:���痎 ��ᜏ���#X�W\�!~1�~�GpߊWQ�&��3��6Q�H���l�~K<G"�^T�;ؾ�׍�Sҧ9׷�֣*����X&�'��1%5?ڍ1�g0`J&�l2p�W�#�3S�1垢�΀)��l�!��H����5�����U�`+0�5�+*��$��-���߲?�\���u�5>���\O~s�)���*�ڸ�a�э���+�8j�B|�������$�f;�+k�����»�ᕪ��k�&��x�E8�����n�S�iâ����[�e�S{TY9��|Ͽ�E/�
�f2i�t�ZB�6��\|����H�_>����Q�V�n��r8x����Uc�Y��'���ܵ�1l��+,��Ii|�ģp�G?���	0��	�׷���W��P���,]n�h�>���
�/�пc�1|���������X����vͲ��H�ZS�VY����[
��-q��w�����?c۠�N�M���k�����=���H����N̙ƿ�X��C�Y�	���C��'�Z3^98X���>q���2p�_7��[��q/�T�dW���z��q�	�9�4���<W]q*��*t�Z�yW�t�[;���*s�5j8jJ2+#�^f��Ê=�+�و?޾/�z#�A�-��kb[^�Dnd+>z���η.�P�ɓ����BP6ْ�=�3w_�?m�KaY�ٛ�}�~������뽨��$2�Ӻ]\��P��m�Aķ���'g�s��������tF�d������ef4ȨVP+Q�	rg�4���Rx_c���^��aJhh����WQ�P+ês�Lɘ�9�\,aD)�u���C�W�k6�
�&TN:���*�<l���H�Xݚ:m�Z�b c&�/�+P�,��C��H���$�����ػ.	�/�0��(��#�ϝ����`�T�����v��o��@���;?����S�_E�5    IDAT�I��+���U��dNn\5��3�q����'-A��s���0r�����N�;��S�t�*<�r|����J�����K�,	s�� 2Y= ��7[�.w�Xr�=�iKu�eI��Pj��lwK�#qk�s��z{�1"f_$�9�I�Ѿ���U�Mv�'m)��={�VƔ�ӹk�U�B�=U��0�,ֲ��?9��ʥ8�����
�6�Xb9�/��*��=O`�so!����Mb)��Y�t�t�?}w������7�t�����ԅY�l.鶸�
�V4�[D@M`�0U�kx�f���H�}f=>�!_f	Ϝޅ���%����b��i��cqUv*ɴ�N�-�@�Bs��=]AM��R�ւ[n��T�zh�%��γ +@Կ�'��<�Z��)�$o��{5`,���y{�X�	�6�bˎa��<��B����)����0���2�M�q�F�P枋3����3l�^�@�g�������[/T��=WEF0�����4���AкDp�D�[4���%8xQ��B�<}���}�)R�p��U�ӽO����!�L�s"�� e3�Z[EԒ�>}�j��A�RPr�[?�nq5PU��ܜ\w7���	X=S����l�.Z��6��/7; U�������z�M��q�	b]�!f�*e�%�
��	�7�?���8hnT����s�����e[�����c�i)H��02ϐ��5p�_^�_�}~d
�F
D�<�X,��O^�o}�\,����;͓M��/�=�F��B�ԙ�twH�bO<�kT��}��܊WZZ#�����$�1�/��s��	L5Wk��륒�k�+/��$<��'S�Kb*��P��"a��1a^��"J�YC`J�V�j�L՘���"�1�|�T��I��*>ʹ<�RY����Hye��%2ZJ�Ԕ����&<c���������q��V)��̘�� ����L9����-�?\v.Y<U�i�«o������(���h�K��s�;5��<	g~�X̚�ɊT� _��P��D6>���X�����7⑧�bp�G$�A*�A�XDn|D���.��T|��S�<�_¶=�7��I�d�)��������S1Z;��"z�G�ڛ��Ɔ-}(zUqZ��˘2)��~ >��#1k�TQ<�r�_�<"��t�S�<�5ك��������rØ�wy�<�=�3���)ݝhϤўII!{���.��""i�l�g)��~L�~<D�>� n�\�v���ww<�|���Qk��a/f�ͪ::`M j�0�Pm;�0�=8{z	����1`H�|i��Z�����[�{XA�]����!L4���o���_/�E��D{�x��	]
C�(�:��P-�e�O_�$��$�o��e.���h���������.�`�cc�9|�*��s;p��g0Q����0&���U��:���yl��:N=~)����0�Lt0�3�o�{ �8֗kD��ڹ�GkA��Ϟ������nl�Q@���;I��й!�j�B}%w����,�]MMh~����A�b<D���,f:���>�KFQ.��1i
�ݓP�G���0`*Re1?��:�K�ͣ�f~3'`�����-��X����Ĩ�*u�9��q1��F�?x�&���9��e�R���"{e�)�Н3�J���4�����Qg_g�^u��>�Z�DBF/�^�FE���uGq��b��0�Lt�QVd,�]B�f[o+�I�s�F�U������P�$�@Rz�q�vMb��PX*U�X<o2N<�@,�;������dc��{! �L���ʢ؟�+T�a��|����[��P4%�cn�lT՜�J̿%!I�/��Iɵ`ɾK�0maT���*�	��
$t,�C����9;獹U�GU n6��-�m-.9����1�⤶P7�K6�@-����5G��^�����b�{��7+���	�(���;3�/�$�q�>hS��RV�=Қ `͆	�#�}u#��I�!����&�u�ϙ��2?�#� !���n��;t���5a�g��9̑�3ԒFs~u�O��L��&���UP��P�M��gQ-��;�I�	t�B�d>/��s�c��tA$�<ݽ��ip���%��v�cX0�����(Z; �
L%>�����Z���	
F��ъK�*�Hq��ʼ��ǯ��W����u�6m�ǫk7�շ6ch��;Pc�-AioB���1A��U}qUR�!�k�Z'�ٖ�Q)F��
��hg�98�4�`O���<W�[Ӄ��J���"B�2��(�d/\~�i8��R�P� ��<��&��H�}�k����Зez5^#��=mN����bJ+�i������m�h�܌��V9d�H+�� |Uq��:e8M=�����Ll)ӥ�q�8���x��M���:�U�7��b@�Z��Rg|� |��'H�X�;�bR�
�ĳo�;Ć-;Q.�����컠G�NX�5�G���?��W��5omG��\�"���¿}�B췠C����	7E9t�#��_F�O�{��
LiV��T)+�/�Z0i-�i[��IX�h�/r�%xi��yy$�`Z�s)�����{�/�G�S���)VPEFr���xU���@7h�|G��Ǥ��\�46!�!*���u�K&�Z<�j��9�|�\�	�^L�i ʩ��<g:�7Wu�+�	^QYѶq���Y���Yה1M���w`J�A�NUw��Y�h<���-6�t�S����ø��{�ֻC�xԜ����(��<�u�p�Aq��'␃�#wĺ[��/�EK���ᵵ����xu�;+`<�nG=�@,���[�b��1a$#�	|��p�e'J�7�N�<�7��I���N ����-���:����eq@ݹ����2�A��
bѐصO�9=SzP��1^![�!����!i4v��̥I���ZƗ�'ШQ��Q��2:"C*Iք��/�T��sX���YP �ek��s�$ʀc���s�L�T����ra�"m���T��b(urU	^�bQ�.8X8�je��#�5���h���
P�b�5=����ǪxŘd��ʱ�O���'�㒦��::�%L�ذ�;G*�B)P(^���,2K\�\�:�Jm�*��g&fN����4�Ik��U=yϤ/8NɘΔauѯp}�5	��͜�z����y2&��ƥ'�Ra����w�`��#dL�H��D����*�;��`����%&˨�C߷:�4�q �Hh`k2S�:�O�*e7]�yׁ�?[pq|�ʿm��|~��bU���N��+p8u�g�bJ@Da�T���h�}9dL�cʱ8gPt�Q���Z�>�����Rʛ��`��~����z�b����1�1`�54&
���r��|�S�Q�!e1����ǰ
�L)����Ř1�`�I�/�@���Ƭ�I��!��)C�ه'�ʇG��H�3K���KSg�<i6��xb:c=9�C!$�qY�J�)	�\=T�Y$cu$c7�@"�xAP��&*.a�U@�X�kS��X��}c���w!N)�i	��Aѷ^Ze5�afZ�QR騏d��TJ�x�bl���5�9�"�b�ϙ�,~�j�9�b��:�*�����S�����Vb��&��7 c���սs���\�؛����8�*N��O�Fݔ���"R{��;�!���a�f�l�9�m8�:1 �K�&��sQ��~t�E>"݈�V>m�R����w5�U�Ye	�U5��)�q=���اGv S�e|�Sq��b
BwY��H�(����_�i9^}�e��\�T�T�������;L�b	�c�d\K�(9��-|��1 � X@*�P����ė�kH�#��E��V�!�s��E�Q�����o�,}�A8���0{�n�����Dd`}�A�h���:5�o��`x��	�{�w:�ӹ߫T��垳Nٯ.�Q}N�?/g��"ѐ��c���<�I��=���3K��s�5�2w�~��<�i��ujkU��V|7�*02��<��^x�?�&��eQi$Јe���&�ї�M��t݋����&����t͖b�
y������Ҳ�@�@,Z�FK�HJ}��<@MUb��懁�0�h�e矊�O:�;����&�(�g8\�X����4vMđ��L�8g(s���qɺ�����Nv&G���);���[�����6���,�*	 ��,+�1��{���r0����cfo��[��Mr+X�����_����<πR��F��H�(�+W^t�|��D�+�j2�"m������o߿ooD��_���#��O=W~�l,���ȱn�~�.#Y�������!�e�D�e|��}q�?_���L2��B��;��Gp�����M�k��,��$9����X��J��q4��x��q��-��l$Im;jQ:>7�G�F�B�h��	�Q��Rj�t�7mL�R0׊9�Y� �s$����l{Ɣ�Յ)�qnѶ4j��1���tC������*S���je5����%�@=u�%���O{��r�p:���Zc��{R�H�)���������U!0��w0���e�⋟:[zL�PK�^{g���>�}w^5�d�èz�Z���ռ�p/��;��X�x�N�F��m�p��[�n��>�w���I���n�����SH$�N�bb�����,�|��q��4ч���}���J�c���##UJ	�#(���JN�J	�V�t�Y�~��liD��rp�B;�4k��� pNZN2����01�WQ�V��_	z�L8��T�(5d�	��_�W±%��#r�0�墥LX#=<\��4�y�8��0��h
�h��/��0G�����J_��֨����|q�Z^z#k��0̔5��!,����q� 椳��AK}��)=|oK6�\!Pdq�Y��M��	#j��5.�:�p\d2:��a�y�(�P��^ɣN���=���Gʦ�GŶ�Z	(B5ks���{i{eiUZ� ����SL �s�D�T�B>O>3	NgQ���y��P=�	L�J�-� K��QAL���y�K��bD,&���7\+�Q�m���ϝcdʬn������0�Ec�
���h>�x�u���C_K��t�UGe_��)O����!+��!��Z�	L��T`�����<4�
�����;'!�5	�dV2��Z��V(#"����=4����=/�ee3tR'�8�L�eN�^j6�M�)%2u�S��T�lĄHA�~hK`��B�+AɏhV�zxd��Zܐ���$�.m�P�� �����Tg��\����d��,��"W!�*��*�=;L����5$�.*�&UQ����[J�Te�R�4�ɾX�7�}�����ޭ���*Ga���دG�$�};Ge<� �A���X�y�d,���$������m{]�o��s�I�� F@��)2W9i%X),'T��X�䄺J5�p}|��{(�D��L�B�%�$�$��3@7j�����������;LB'�������g��!zY�
l�S��-͆N	 =��  ���j*-g�5ׇc��o}�<,���'Ӥq,R����V?~~��?K�4�PJ��Ϟ��et��&k��痑1<?�8�m2_�t:9��Y����ɀ;�� V������p��Z����8��"&�E�������; ���DW��:3�6 �,&H_����~+�9M��?{>gxs�p�b�2��L��qݲa���a|��r�*Iuţ��\ݢ%�@�k-ѽ���A�(FOw'f�5ӦL¤�,�3S&w��#�����6���Z�ZM����P���O�qGSe�ٿ�i'p��O�ѧVc�P�*qF��M�	�"f���H�29#�������r��熪[V�%cC-��g��)j���~ɹ���7R�͹���^x�~t�+����8ӻ!ću�r&,#����|�>�&�$|�6���-�S
�6��3�I�i
}-?���X��\�N*�*UwE&驶Zb�(�Y�+���*m�18�J2��Z�$jU̠�����Ƴ�
��?������l)x��Ha_��,|��}���o����q�����?�FJQT�f��x�hg�t.?�,�Ӯʦ7��f���p��/ⷿ ;{GĄ�C���$��b��'0�	���!�~���W��2k�&wIa�J�
��|f�����3�/*+$�g��	������8�0���U���/ZWP�9��"'���H������I��+�^h6���d��\�� S^K��C�@���E8�O��k��f��Y�� �/�F`�,"�Tӥx���,䔶ui�K�̔��e�RD���Q\y�	�ܙ��g)�רsr�(���ݸ����)�ȃ)0�w��y o���n�k��Z�l�N]��>5*W�hx��E��Y�%#�ܝ�>�ajO�0|L��F�104���,F�x��񴸝*�J!M 'c����rè��Y��U��8^*o/���=�n��	���2H���P<�@qb��aT��z�I�ę�:-�+S�Dl�
���H�u#�PA:cɨ�>:�COh�6D73A{�8�D�\�^E�S$a��"�L"ݖ	\V)��Æ�E�,na7�}�5��Yr��EL�T�[�%��uL8y�S�H�@W*�d4����Ǎ�_L��(�*]_M6���c�Z)$�t=L�`;]վ"�!$��OP&�g�e㈥ۅyc�;�JJb)2gI8�h��@�^@Z�WP*�e�Lq��^.	SG��kKfR"[l�8p��U��))�=~��%������ �L)%�+�iC�M�VQkVҘ�jH�#���B1;��W@�S�����|9(Y��uarEc$pdE����e7��K��D�B�p'BF�M�^�Db)�8 �R+2��hi?���sJ��� �!�v��!�<SV���C!=�Rɴ�[B:0��^*�0�=�#�9I���x>g{��D�,�E�0���"�%0�����+Q�ڞ.ԓ1��ŤA�c*{��\�o"���q1���_�8������v��Pqc����c�u��钁�&���5��T�T�>�8��I��rl����f���1�J�d�l�&\�[H�&��b�c��>�]͊��qaإ�!}`M#�g2ۅk,*��V��]>�J��Ĩ�`ϋ����ڬ'�΁�rUdVu�	�8��Ǩ�;5�T���F�9U�]�dʹ&J�Yx1�
���05Vӱ����+a�l���ǝ��jIP\/d`�d��e8���$2���〡�3'��d�1�P>�S�A��a�$�8ʽ�k���>K�m�d_��}���z(���q�ы�ϟ�Y4�4E {��v`�������WcKQ���P�R&�RH3 ��Ne���*\�&ɘ��7�^�J��f967���f=q:�\�
��N��n+%����4���۱d�T�l1>x��0gv'�S�K�#�Z; Gz�䵭��р�4�58�cˎl�1��;��w }����(����YTT�JGd��ewu�jAR��Ha�^�1�KU�OgN��f�l�(0���v��0{��5s*fM���{M��930k�L�˔�r^�����5��|_���pH��	`��A<��Z<��kX�y~�Ɏ��%���0�پH��B�U6����*RG1g�VF]6L3�?:����[����L�l��9ǜ���/=ԥ�0��at�j�����ׂ�
��T�PEy�>�?����\��p�f��F�⩅u{���}i,p1�$}v˕�ҷ<�g��05�>�ٖb�ko��nz]VM�.�?s�������>s��l�N���O�{�mZV�����k3��;U�
(��DDEc�ƚ����Ę��9'�^�[4�Ē�����("ED:0�+o������y�o<����g��{��y����^{���`���o��
��m/å���y�oM�G>>�W`mD��E���SԊ�sm�w��x�.�a���L�|M��&!�n>����_�۷�������a�    IDAT���I��"���9y�����/|�F�ful>�046-bD�cG����r6�ƙ�8�y�SWZ}Og2�%{sqA�b4�%����t&PX�U����T"[b"��i�$W��dV��(f�r/�cZ,�eF�)�)�-��cJ��S+�g;�꘲�<�?����y��՚4��"0fԥ5.��a6���|�p;��Qw�/k\���$l��4������+�R{D`���]�S��[��T�_ܿ���e���'���D������r���ꎀ@u��l2B��I%�a���y�H��93�*�f�R0���r��Vk�]��H�Y�;�b��e�\L�q���Ч����Υ���ܴX�a�/a�ReU�F(��B<�������{�RS3+���&hrX��ʜ�3���>y��3o�ClXn��	����D��9��0d�=	J���YE}�c�6�sv��x�;ZJn�*x(t��w�P�챃E - �7�L�|G�<�U��뀟H'Iz
�;�&T&��=I"@`ҭ��L����Uw�iTԓ��?u���*RE�ڄP�2����r2a���bУS���F�e`"�D@���粲�`��~����%��8"� �hn�!�F{4��ȁ�m=����WQ(Tto�5ͳ\.�pb�Y���Y((2@=�Y�B��s�ɐ4����\=%�8�:1B�N:��x��.�n�m�-K��u��s�qݔe�C�U��%͓%��`�Ϊ@��,M]S"I��`0��(☦��0�B��&\s��ޒ��*/�׽.��wb$`����F9�٭aaD?��e�376`Z�1[kc���
�ܒ��o%0����Mp�.��wU|!�N1^� ��+p+�
,�]3����Ut�̱֊@�u����N{�m9�Ә��j���� r
���l9�ڍ�V��h��1u�3�ި۽��K��D=�}���]t}F�צ�vx�꾪�n�����gK�Q����>;)p:$�d��C���;"���1`�T�@`<�`�`�b�C63�{�6���Fg�w%Q��k���E��,U��x:�Z5�W�PO~#&� ����UTt�t���iB/�+��Q��q�	rt&B����3N&�ٳ#kƘCթej]�H�è�(�� �}I�i��o�G(� Ҙ��ώ=�鸵<�����ѐ�G��[wѰ��[�/_���f�E����L�uZT%�E�7TB�ϓ�6�,��N��V�Pܗ��i�.H�"�0,��<c�K�-'sjy�F��X+�E瞎�ؠ�rs61�^�)n�|�e ~O��b���{h��a������G�Ď�:#tX���^
I,�ۧ:����>�T��fJ�&�A̖�;`��)��#>�R��&�<Wx&�w��z���rc��JXhT���9u��8�q���a�"j�!H:�^�aT��?�����)@��=��ko��?�ۖ����0-�e�4fn�3_�JX}{��W�Ȋ�ٳ�Z�F=Ny�Y=tܩ���kꔪgqN�fJ�:'�8�v��.l����g?��;/���W�����:�������ǿ|VGML�岔�Ġ7��47q-	����-0��ĊF���~>:�Vx!0�����zPj7��8{~�%?�=�)����+xN���8����~E��Q�� ��Et�,��/�����C1O�OR�3��}���ԗ��ڨ���^�c����¬�Q��E�?o}�8d��h�>�ï�s���;�?����ʗ/�Yg>���N<>@;���2�wp`:�c�Gc�s5Y@��%�M�3t� t�O����`D*�Q[Zĸ�G�9��E�r��+h���HT������)?��5�	L�e˗�cyH)�G�TD�)G���j[S��L�\yz0�����P&���M_���u�:�WK*D�\�&�b�M���h��8L+�4��������_��/�V��^�S�!0���<�|`�����m��wj
pZ���:�m��y��#�|=�}X�!`���Q��t��A�O;f�4|1�r�<cW��B�v��eTrk��7�����r��W.�%��߮�ε���F/T�3s����7�'����U\�G
�-X͢U�EN��M��|p�}�����L��Δ �U�YU�r,�$�R�n� "J�L�9�dF#�5a׮]�d�,Щ�b�L�E`p�JD{�Y��$$z����+z�X:U4�x����	�-�E�%����%���������4h�e�3D��ɜ2��_�iX`�� �X�S:�2��u�^YS�%�Ι���\�ǵh*�����R�����9R?+E�9�y�2���	�]cɟ�D���� E��u�X%r�X��+�<�2���;^�h�Nn��bT���(������5�$�ijk�VKP�ٓ���3�a�='��n;e�bA-U�u�y��8QJ����S��E\�c�����n2ù���EQ���x��'���4�2g<ĤۖƔU��:�1����3S �>����@�Z���6+��$�6K3vL7-`)��Eg�q"��{Er2Cq4SǴ����Ui�nz7uK�S��,EV�4U�#Ir]�[���{��$�:�íc�$�AOf��$���@�٬��j�Z��	Y��qmX2�������� �~��4��Ll����F��ɵ&�(׮wPyr����a�R�^����QN�c�n�ę:���vO��N�,@���0ҁ#r�.3�.	he�G�=��g����ѡt*/����N��NZ*�/a���w!M�8�\	��G���p�Bۦ�ā����]�}.¾�f�Aȍ��`�$\��[���C����|x~���A��x���Nm���4����f���;��z�����.�ɇ�t���� W\{>��o����%�WT������_�r!����|�{��i�Z*Ɛ�[����<�X�bB]T�
�,.�Q���+7ZþJx�ӏ���<Oٲ���4P�m{W�ҝ�y���2<����k3<��N��������C�lC��s(/3/j,�A�q�0Y1�EKϑ��|c�{�8�Ay��o��{~��`�v]��3�����V�"��óHZ�Q��*0h�y9?R��#�s�u*N{�������g@��f,6�����%���ȓ#|���q�U���0*,`Rj���d��>E�	�X�RA�5�>(�j��ʫ�"��{�D���:�Ө�q"����-��Y']���q�|���o�q�/1��V����}��_�_��v�1�i��.3 P�=��=���L;mQ�2��w�tw����f�����5�19���Ȩ�͜W.�'\19��e4�ajg�H�L�@\��	�ʫ�X�����K����y�����S�_�M��;�Ǩ�������]��N{;Q���g�����"<����]Խ5�t��ܻ����!�7��"y��b�0|2�޶��\�qe�ICT���L���T��/&�-��G�@� ͣH�b�ws�E����"&�z�{A]�Q��=�ID�`JPOɡ��1��f�l�I�χ�1,�،��0�tLǬ�Qf6���Ya�іC�n!�T^�\d�~��aܥ3����d0RTy����瞣;���P�g�fey�Fs�����yxӅ�I�t2�����G����:�g�p������i9��6���+p�/��pH׵:*���Z+s�c�X$�T�D�V��D7$M��	��iHʲ�73�
ux�2&�!�V�a<ZF=��;�|1^��S�1�n���^q>�k��]@�?@���f#���w��UxʖF"�8�lZ%�Ie�*c��lk߸����~���;�L����5	z~���4��bXg�:p�;L�h�N:/3��mѦ��\�u�Ffb�:��q&�\�4a�+��EP+�SjE�t:��5o�3�8�ٗ�)Y������J�ڳ}ih;�eQ�����L����W�G�f��*���B��[-�Ҡk,�us}Ys�����@]瘭)�)$��z��.z�1z�.��6��t���m�ڱ�.�PZ����ʴ{TM��nt�h$cZ%��[^gIV�*$/��y9UѿfT�9ׅ�Q��_w���Oͽ5*����1nt�M�:�D>���v�>����N��zUW@*�M�^�ć�k�� $���ّO`���>���f՟��-i��w�xj~i�iL+�1-�,S?�h~�N'�3�!͏Z��н.�Zi����3�ZSG):�4"�1^�Ȏ��;�~� ���p��������R�d�{~=��QI��?�(+\�ӝ��y$�[��S7�P�Qp�/4S�n4�~�ޚ�*���߮�]ӯ�� �����k�*���T�;�^@R\�$_�_�l�(�Īu<�-�ɑw�5<\ �5��5L1����ȟ�PPO	�7���c~�'�Rb��n[WD��%�r�d.��k>�)�:ƻx���tU����7�$��	��Aa���Ւ�l�z� ���
�����u(�.�S\-	���~�geA��?��X����ʦ��sS��}��w��Z�mط�Å�=�~�����.n�������E�&����	-)1��D2+��&sܯ����,�:�H�g��5��Tq�:��{*�0��I�ǿ�X[ކqw76�p�ӎ«.y>N:z�F�1w ��h���b����ص<��v<��x��m���{����ع��hFS<�)j(�t]C�R�X#@�	V����e�=�9���0x��|x7����E�S�(χHl��f� +�q�3����lP�54O�~���-`���*�v�Q8�cq��[p��b�MU����h�[duY\��A���_�~���� ������+���v�<���J\蒝f\\+Zb.y!*�FU�=k&�a���EKYR f�����v��iR^�c&�F�e�-���s������ݹ{�������xb�EU��Y��i����������|�"SV���g�ˉ� ����d��-��u�K�bY&��?�1b��B�k|Yhc3�[�7-�c��9L�y�8�Stfm�QXƟ���x��Ĝ?%]c�L����m���Awf�t�ܯV��A����2ʳ��U\�S��\�#�o8��xl1� �޳U�O;h�*6��Ɖ���>����o@oR���F���
}2ؠ���G��ktt����=��zW�o�X�~��]T,���&���,d77���3�p>�cJ-=Ls��ϪU�瑫W=.���;�C��/��.�1��p�l�f#���\��C����U��\i���$��T��JU�z�]Rs�O�����Y��{uKLgJ`Z�t07Y�[LOĆ��=�gn:��(��Rc�N�'����b�z��
�w=�V���_mG�OÞF�٤!��L�f�ܠ��Z9\�2���w�jn靦s���Vn	vj�gW*2a�vvc:^F���;�|^z��l����~��_�c����h�nw��������W�c�w4�DM0����HB&�x ����o�
�����א+��i ����uݮ��vPmvvۘ�R̥g�h8�� *�jI`Z`��!n~R=G4�!`�&0V��������O7�59��2hx��ڇx�:�k�#����-I|T�$��d͓>ui��o�����1��Gf�2���4�p�jk� �rA�U�*;~cQY��	v��.���V&�t$���τ�������f7漏)�Y��®����b��+�Qd=�^	gOz�*q��LE�A�D�!��T^�d��k ���:l���b�O*�\�!�a�Iy�r��&%=I���$��ɒ���[���1z��~�%k-E%�{tLsL�15�#&aRL~"�']�s�f}Ryw	�6�P[XS�#v֨G������V����X31?L�-v��(n���t 7V��1ʳ��n�"��p��j���qG[����v�������B9]�����:�n>���*u##9�,�
C�	k�Rq��xd�U{na^{��	���X�F	���_���|�,�(X�6s'��!e��X�A���$[|}s�!ܨ�y�R��(���:|vR��j�8��F]R�����e��D��t���`#(�����|�n��"kOy�j�S��,.j�j?�1o���w�"q�Ρ(�I����=�1��0I��ze9�n���15�X���4�n����w
����6��L$Kl���'ۑ���Y"����6�1���Q�A�%%�~���V�(�9����I����yAƋQk����FeLK�0	4��?���W>���g���l�*�8�}�dx<�K:l��;q�~M�����眆��-��J��0y�����Љ���3�򾭸���q�]��'v�K#5�WJU�;�a<�I�a��+&��\��x�u	��(����J�����%��%�P-4Ύ���.��l	�u6���QC�EY�vQ�=�:k�5�0���m�sc�y'{�w��8�ԓp�~�K@���v�LZd1�m;�$Qwܵ���������ʠ�ꘕ8Ԝ�)�J�t>B϶�DEQ�6(F���4�����}I,�����)�$�R�Pˎ1��0��]�����1��{��{/��]�X��Ĕ�Ӝ�Ji��u�����o3��>Y`�]��v��ʝ0*���)�󈒉�yg�����K��v��o�͂�.�F�Pk��5+�[A�U�G�&�v�ӹ�*��/���=�p��|d;��?��uV��+M�IIm4�52F���ܤ��pYU>�T���}�2"[Sw\]\���RT��G+rI��n��J�θ�����R�R�|2�()�b��y�&��rg�8�&
�I��$�m岀)��}>7J�
�(j��tv:r�e�(ј�ѿVCqaAS:�X|Sa��Ry��<�<[[]���P$Şs��uQyi�$*�K�|��3T�L�^��ðC`:P��4��K���,��\F���#q�s����FC�F-�M��K���^r"�(q[��)<]L��1jL�����୯�XT^�0M~�p��W�;�@@҆u�B��α�|Q�lu���:��]�����#��I�q��1'BT^Ҁ{�F�����\������1t��d�P�8�a�Y�a��-�~!N=i��@�L_�1ʆ��a�|�,0�-���\v�q���Q�ؘ������J=�u�`�~�~Q%}f����&��qx/��D�}�ƿ�k.�ِH�2�:�_n��t_<S�ǵZ��2`�(�h��9oJI�^�*���#�$Y�J�-B���w���W���%?<	y}i7�U׭%��}��/��}*-A��vQ�r��cJ�1QA���v�Q�"8"ՁI}��PǴ1� ���+�W5�GzZ�lu�݇n�
wE�K��08Mc��W�A��b/R�=L�����{��Z�ـb k� ��*�t	z^L�^�����+{o5�\��p8���@ɨ+�fZ�@bf`���HXH������h�B	C4�/��|}م�1�-�n�֜G}q#f�����''g�Ｙ�Rx�q1kU c\ߛԔ�^�?��C��U:m���qF1nǭ��2j�G��:YQM�=��TRϺ���t]��,	�!ǹ�d6�g3r��e�$�7��w�h �7�?.g����T�i�B���E�	J|Ҙ%[�Fa+��ޚ4�~�kT@�>�a@]��n&�"�Ϸu*"���ɗ3'�M�G��|����nr<����`5c��l��t�V�r��'�b���U�%�qf_y���eI��&z�*���� :���.UP�d��`t��������g�X6�ӷuH�-E�8C,mԊ��%��"3�^�į3���8�}3�$A�K���H��!��ї��J�7[��4������ZT`"�!����%eTH-����>�w�1N4�
�#�xF�ڀ��X�(��G���⸾9-��n�t�����";%�.&�>ƽ5t׶������W��y8��&8>%�w�����]v�����;qݍ���{���]��֤�"��:מ`��/�q/�#��(��$y�ӭ\���$�a��(Z$���{'�%�<S���Ue-9/Α񣈨zTPC�k��%��n5�a�gO^~=    IDAT���ɠ�����8`�%�q�	����ḣ���hb���RX,@H��f���?x����qϣ+�i��̂�	�԰3�����W��jy=�oz��ʊ���f?|�F."֑3Ң0c��E��}H��������9ӿ�����z�,��/=�#����$>	��@�Bc�pJ�+�8i�	W�Xi�43�)�"^ع�yv^�q�)Ϥ��qo�e#��N���pT��5[/�Q�/�^�"���GaQ�v�d��hO�|����_�ay#��9��Qo�]#)oc2XE~���\�s:�����EuN��	[���f�gx�T��_n�GӺ�֗�����>k̐�o��o�J�5�e���s�|��q�����9!�T^��RrįE#Zg-��eʤ�v�,�ah25yj����wV 8@ǿ)cL#%g"ZHͣD�#GF1X�H�D����L�U�K��x'��K�HSg���s��C��Ƙ��ȡ\o�P��a�tg弶��3Ћ��1�y����P�ba��?x�yx݋��"���O�t2��H��5���_��qP(��'�����S���ݏt���?��Q���Q�����R%�D��e2�5�l'@O�����&UY�w��X�����Ml8/u2څ�j�G��K�;Y�o.^:{]�����O]��w�8��>ʥ)��1N:z_v��橍e�:�h�G�Q����?
�745�A ������Ʒ�tFU�Ks(��a7�	��`�C"���:�2��<�X�R��r�I�ʐ�ҨNU\�VUNA��G��j*o�u�`�N��Q�y1��V�.�<���&K�|��TK�M���Tc��w��0_�ׂ�oЩ(�Fr5-��ĖJ���s2�*�%����z];�X)6wS{ 6��V<@�^��u�%}���~���](��w��|nQj@ĺgI�iIEҥ�lP�%�6GLO>�~d~*��'4� ��݌����B���Q�|�p��N����B�D�7�[�.����lYס�h4^�I��y,ұpYX�Ϧ�5���t�Q�������%T��L��L�)�7���=��r(�(1��4�L��Lp�su�6�cZĀ�F�8ꖈ�dN�}y��ѕ�?FQs*�XΡ��&ݷЌ�d���
�`PC�i�J�CL<�!�K�th� A��i���sP�!ku뙨Ǹ�0�(~�H�"Nm:�jr�+V��g1����r�ގz2����.�����o��0�g���֙��D��R�Az�*�S3a3�7?��a,h`E2�8��!����/&Pa���K% �d�'����0�i�&�d�h$����0a;�q&�� �����K�~F���K�s:s1X$f3�W-Mߏε3�DJ_M:��Z�Nr���S=Ѵ�2 -fD �����4鰹�]��N�k���|��MĘ0SIϊ���q�ޑ��G�P�M���D�4 f��P^�,�eq��x�q��nk'�+�t�~x�%�✳�����F#J��%����7|���|W]���{�f�s9�gE;e�=
��c�yyFQ4:�V0鋞yRlN;Yq�b]��N�b#-�9��'��P��*ȸ�*Ċ�HF��h�>E#�<�P!�a$ϐa���U�GO��o��=�׀SN܂��,�uƉ�w����,��P?E2�'Ied�j��KW܊�\~��Ŭȳ�!�i�T��+d�⦆���ǞeVg�{n�~r9�%bi��׶���vE�Od�ȭ<����V��v�,q��5RxfnK"�
�[xH�h9�7FQ����I����U�����Z���貅�=]$��l��Wb��#
�62�	Z٬��(�_�$���ʌ˴�f�9Aq�Cy�o��������h&n����Ż��SX�-����\Q�x�����"h�хC2'{�QE�y"���q��5���N@�k.���l�;�������vz����T��Rʀ�%H�������1�(b��չ�V�,�U�(Pr�L�"���^T�<���1�r\c S/�3�T*(,�il�8�ǐc���G�Q�X@�TD�9�"�/�&P�L�6n�1.��eq_R�����I��~��~��⛀)GưX�`y 2������Z��%�>J�5,a�|݋4�c�b���uʱ�`���~����EW}�	G��o��8n%�Ry�����
?�}+��2���CwuH���7��k�9�bׇu�0ٛ���t?�!��&W��4W�v��.�D�m���z���L��?����x�?OTi�OJϴLژv�c�aR��Y��OG�ժ8zˡ��w�)~뙧��˛���߽��p�c]��٦MTȵ�+���Ӄ��R#E��C#5���$�a4:�����T���k	NM?�	���3�a�f:��
��6AY�P��2N��F�w��`����9\I(���x�S�&�#���~~�� 0}׻����=��6Wb;���H�)�ijc+�
�,x���f0�ۜ�3]��`$pD�)�
���(z���Qfc-Z�ْb;0�G��מT^3����eAhT-M�l�J��\*�z�4p��V����x��'�6��t��|x�4���8��e��y�EQ���ҢS�WA��r�S%δ�E�80����\Du~�We~4+��SĺVIL�i�����6W��i�A�`�]aU�`Z0`ʎ)�v(���2n�|Ҙ�L�$�FG�)K~@�7X@� xBE1[X;l�Ot��Ź��Kg�nhXx-cg��t����@Txl9�Nih�v�������:)��E�?���֚��|b�6*�����N��'��O,��0;��ŽF �QD��D�U��T�Zf7b�%�s9z�pD#.�f�ഀZ��3]r6r��K f�����+qR��WO�b����+��m�l$��(���[�/)��y�[>� �|��(�a��!�7J�m��5���8���a�)�ţt�k_%��x��b]e�~>S�Nt/VE܍�j6�W��cW��$YqgkKԍ��ڍ?/�=�hg5���TA39����e2�M�o�#��qM�P��ag��n�m컱�K.x��)8�������%יbc5iۗ'��-w���݄;�݊���\�n�,�ѷ��]ll �L����(�����Y`E��x�̈i'+�	�̙8{��-_�W����ޒ�p4�3�2�E�O�	k4�%��F��"#G���r2�c�Y�l�Fn�*������>�s&޿n]Ԅuj�����J2ݮ��I|���_<�ָ���

�\f�'2�
g)�*��u�Y���2�%4�����79�z�2��2�d�M�9��߼Isŋ���=�~�j�$gw�;�L��3��z*�,�ؿ^N���uk"�nR`����Cq��Ncp
L�!��D:ᮼ��Yc���*�(�q�����x6��[y���HO�������܌�q�|3Έ��RI���z���Y~�B/<�d��^���*����u��$˜1�����L��?mb�C}q��,R��Z ��ʊ���^�Yq���.׉�N�&,L醫)
��u���<*ә�);���r��
���T�J�yja���~~v��+
������T:�Y����I��1G�80�y"��J�P��	�ҸHƩr�!f�)s�p��؋��S�<���{f�Cy���U�����?�e�z����>�e|��Wk���O�"`z�S����{�c=|��W����hl�4��1�0�T^�NZt>4Y· k#]8�S��<i�|�oRA�a��Nh�6��e�&˨[��?{^|�	Ҙ�� W^�0��cW��cng2������Ơ���*r�.�cz���a��������/x�fxqA���ß�_��n<�� (ΣXn*�mh�x
\š,�fX9X �K��)����l�Y���'i�q/�1	c�8�#�U1y]w����Y&�Yn��H<��u��� �1+~�T��4,6�*�x����k� Ҍe�r����0I��W���e`��לU��{�0�t�s_YU%-��V�e������5}����������<�ͺ*��)2ך��'̩����ޅu�T��H�.v�A��ۙ$�l�������K�T��`ѯ�����c�Jw�:��W�ŋ.X����M�&-�����A�SF�����s9�*�)�2�Kg�'�Ś�Pa:�Ё)��4�����	�J�@��'�|���e;������ɬiL�(ScZ)������b�-�+Y�����VW��
~&�i�L�D/��b�kb���R�����G��Ta�"#i⬂Vkh.,�`,�iZ�{l��Qk��ڨ��2v�8Ì��k�Ù�c���g#���aۣd���1#2���F4]R�XXܠ�R3�:o�:8�ْ(u�|�dd���LJG�2�	i@�AEc~^]]�t1
�� 5�'r.�f2P)��A��L>չ���Q|M�(����ݒà�G�0@�%��ب׋�n`H�l����E�k�Ew�|��W����1sH�44��(�Y+n�fL�b𘝤����4���Lpi���Z��	���v����4��/<�wIP��M����b�z)/ѨYq�.$�u�"[�7�Sqߓ��`,��?����3I��;�]~U�����k_q>�:�(,qުˊ�ȠQ�����R��Xn��=���;p�]�`���a���.����r���k�՗~� ����w����(�d4��|�#�v��){@����]~.`ʘ�����4���U�ɑ��Y�gpT\R��3����mZ�1l���fg�����3���:�˺L*T�~�,X �����7݅��:���NL�(V���P*P�qzQ��Ga&ƟX������k|$/y�U�-��/�d��`Q��*@.�'���S��(BXv��j�u���}8�����1T��y��{SL��}���w}�$.eP��RC�)jȂ+l��ً/Z�d�x��,R�s�
�6٫����7ᄃ���Ţ��F�p�js��-���~�vL0,-`Z�)�`nH�7g�k�Q��՝�c�ىڬ��y�s𻗞�é!wp*�Z4����A���C�a߃�@�Q����e�/�m�`��Jb��;]���'���5��RFmÒ���h��nZ�f!���	L�}���T�*�i�#jU�8�Z6?�t�)F7�0E�#��:�ܷ�
����`T�its(iT���t��c:��t�U�M	f�Z����tj*�5N�@�$�W��6�W�_��b\z�Q�ؠ�z��R�c����SRyO8o�]��QΙ��=[��৮�<�ᨄJuΌ��$�,�A��^�XnVv�82@�[�J�4`9�2�s�Y�
�f��6C�E!�0YF����xכ��g+`��Aq��?|������M��v;(䆨�G8h�*=pQfH����]h�W�h6p҉�����c�zvri������>t5�*��V �v�49n��T�Bc!8�z\��gq�=�U �/S�cfG��d<ׄ�άjcfa)�C�ăN�R�]�������FI6GN|~.Z ;zs@��3Sb�8/��:7�%s3��o�Rm�H𜞢��3���
� �x���Me.���M�5��9�3L��*�Q1�ȳ�@)��7�Мob<���ȑ�  4�~W�Ҩi�a�u���;��6�Rʮ:�N�#� U�6�{\W�Ֆ��d.5�P��PI��qٸg�&��,0���u'�Tx�C4jLّ.�S`�}�IX\w�j����k�.����Z}���su�XL)]�`ץq1�Rgʪ߮5�VVU���ʦ�� �qP05�fa0�h��B�<>��T�u]g��w�|�X��"��fƎ�2�U�����ݝ���U*��7���\؈rm��2ر�&�rhG�,��+��WѬN��,a����2���ͺ�Ut�]Y^�Z�-]��,�&r���GXmw���cy��ō��=����D{W���ҋG\Q��w�C~�G��G�T���g�)*ͺ��4������)��#9�4�gV�8�e:%uTkM%�\;ʁ�0K��w9!G�?�:�`��i�+�"<f�s�t���p�����4�����&��c&�Jb }�3M����@����\0���<��G�P�]����7�~��\��Y��W�U�ǀ'k�'��5J�!|K��)�'��j�A�.q
��I�+��"+�46@��,cV��9���e/~6ٯ��2�U������D�E�V�����~����5�W'N)י�$Wƀ1�n��Q��!TT5�V��0Ș��Zٖ�5u�\Cq89��z�bZ�˜ju��fO!yx�1K;�� -��Bݹ������B��N���]�L��6����F��:+��0�-�0��S�ū_~>N>�@�{y�4�������!��3~�����p�-�=�`R�C��gB_J}��cZ���(�f�@o d�\+|�)��� �i��o��0f��{�B]�`�8��3E�L��
[���z釤UN�4_�(zǅd���Y(w�B�� ��+7v���1�[c��ݟ��ͥ��(�&��49�L�;(�(O�q����/~��8bsI@L�{�j��� ���5|���<��q�JӀ<�b�t~�)���kOb���K_�,��/Ė���sVj��_�$�#0���}_��'��2Z�y�i7�f&m�X�!+tyZ����v�9�Ʌ7k~�8$�5���D8���0��6�� ���zM�T��M I����GvL�l���[��sgr�i~ğ/cBp_XO��$��c����Sy�1��*��3/͏�OU<H|�8=>�\����ѡԦ-lȯ࿾�"\�#���(���g�/�_���SO:
o{��8���dx0@�n�����.~���1S�=g��dvd`L�7v���"}��bd4�����68�]c��i��v��>�8Y4֠C+�U�T�J�o��s�iL����m��?z}b�餀���(�8��y�?�x�|�A6�����T�O�,�T" �ˮ�d��έ�?�J���_�;$(5��{b.��]�>`C���6��f�3^��V�3ʻT,�]�9HԘZ(9� �����ڦ	�>�8�̪�Z�Vc#9�C4*ݩ�G�)�u��H����h֬Sj<Ǔ:4Y0�6��q������`4V\�M��3�?g3�lH�];�p�\A�f;>�����옚cY����8���h�ިc<��嬲��: ¬ȫݺ�����9�uvң�s*��|$���I�%˶��Zd�7�`�H�s��;���H ]���GҴ54�VH�5`�/5�J)��X���<�V\�$�usR�hh��i�Z�ޔz
�����X&�,�W�۽��p$`Z��G����,
O�⽭c
��v����#�t�m� �����K��agb��Š;�a��8"�3�O��2��S���~��l�E��j)��e��-�T�~����X��aaqNT[���rXm4��W�?��]AwH�C�&i�"]�7�	�Y��֓8��M����q��b����=M>�uƏ�e�+M�
G�J{��ݎ���9�{ͭ����4^�~s��b�8^�������.8�4u�~h֪ڋ��@��%t�e�(���зK�4딜e:�a�J7�z?���><�d�
GF��/��]ʭ����"k��c�Ҹ�ԡРy�U��w�C:��Z&	���إ�=%k�c���T#.�I��� �����Hdw�:3�L'�>#+��^�qb��ps�|=�h�L�{R��w{P�V��6�.zL��Й1�-~��mR� ��$�@��]f�L ŏp ��^��bG2ۨÌK4��ڢ�M�;�X㌓�.='�A��@��hR@ftA��_?9��~q?~p�����c�7�4_�d�d���.��L��j�M�{�n�:A�̆&�n:�I��&)��CnfHt���i���ā5����]��I�Q��$
0.�	���.g^�ե�3�p�Q8c�0��X�Q�O<KnƢܘN�-L�-�"ol�q�YOǋ�9'} 6P���7�t���D��P�t��]� ���kR�    IDAT����5�+7�/�p@�gw��:M��3����M�y}]:���z�>P�5����E����S�e��E!��@J�.�^/�{/�E�Q��g���C�^.-
��4&��t���I�y�D�htF{��М&##��mj�:cd�kH�+y��ҋj/�H{҆�'kh���g��w��B����)YG�"`�e˛����n�o��^�v����IGx����]�nǤ�Utp�o��w��exʡse:gcm���5��2����:�t�O0�5��![Pkr���ZA�9R�bObu�\G��n�x����ݨ˘/oX2VXtL�b�,�Wf9ԙ����i�cJPgw���f��tܲI��>�1�!,�V˚��N]θZ�q1�fr-aZ�Uc�� ��f���hJW�vg�7_q���L�u{]��M�d��3c��"?�<Z���*��-/�K~�04��N�	0�Ǐ|Y��PN��i��+`��s�>������p�O��`TD�����r�>�n��㤗G[�"/_$.�E4M�/�T��<,���D��B!�a�+�)��\����yg��������>r9���lVB���Ji�c�܈���7�-U!���I�AiO��/o?��*>����W����ghkY�Ȍ����2
ܬe�jn(��h�>�C:����J]m	%���ۣiL��&*��x:����q7A2�݅l���{A�
FPM\���D��@i�9ѨK6��;������jV!��Apv*�+͕2:�:���jjFZr�� 4�%�C�a�{�zaG&��A���3��;0��o~qA�-L�:�6�J�'�[N�j���+�#6�k��FBa�ӝ�3c,�Zb�����%�Q,����R+��h[��A�w���&M_L&ԝ��%3=��H����O/K�<�#ݕ�R�G����KKaɅ�xR�	�'#�Lw˰���:7�|��V����0�d�Þ��;Yn�����L�I#&����#gR`J���t�+��'�������)5��&�Ɣ�sE�#��Iխ��B�t䌱5~�^r������~j H�./���-O=.���6�eW߂�]���VQ.Q����2)�z��Vp�o��W��i��ј >��{�Y����c�J�IZC���[�o���>���Z�DR&Ɵ'�㈐	J4y���^5��5�g�f�?�������&7D���2��9`��	��v���q3���[1�Ձ�iM9�&4���L�?���]Xo*d�e���д��/�C} W,&�&��[~��$6:8�avLM�P2%@�O��'�h$j��g[W�
�Lti�>@L|/�8���K��i�)Id���f�4~;��b:BI4c|f�N�!LWj�K��14ܬ��)��G��){}�Wv������>p	�s*.<�TyP5�O�R��S:v����~?�s�͸��G���5�M�~Ṯ'���XO��>>'��F�i?~���*���HFgqt�p�����U�+d�����x/�[��
r�}[Z�t�zo���۾��1�Q�0�N�L�����hf�̨�揚k:�&�����Vw`�݅#��ǋ�{:^��Sq�a�`��IϏ�^�[k�3���wu��o�W\sF�9L9�Z�,_VQ�#c�{L�sω�H�s���Z��"��/�B{/�����eK�s�
4��zRPS�ᣃ�g�o�f�ϼ新���Y��s˺��Fl����v�w�5�y�<{aG��aGТ�e�$�6��0`r2��1f��$t��^�	^w��x�gc����g��e�_�1����(�6���+/���qw��� �>�T�0hm�|e��������C���n!�e+]y?�]|鲟�7��C��Hcvg5U�țvU�ﳌ)������x?|�Jc����h� ������������1�n�'A�`:kpdu�6&P�Z�֨�WK�Ѵ��AwySI}�r�g�tV+cV)��@:��s�<O4¼�����l�4���H����ƒ��W�\q�s�����T'�ث���|��q�3C��Lc���1�~�cǴX�)')W�ӎ���MEܷu��j�(�im��d����`2D��*zGE��f�VJ�`���p�^�B�cWj��9pqє+eQe���C����=��V�!?]�b����[p޳�Ѣ�sf�����?�<������W������;��+nk�!٨$6nA�EQݒk�P�?����}�f���Ǥ3�ŀ�9ֱ�3�s�;	�7*
�2'�;K~8�D#�i1�yv~�Zȍb0o?xe� .��RÌ�nZ�m��d�9����ц<O�v��n}E���fE씲�#P,�+$h^;i�)ڝ.Z�S����!N�������c^"�-�Z+�F�%3[�U�"i�}n�h8��ʪ�eP��`��6�`2QǴ>�Ħ��B���:�t�4�tܷnlB9�tA��7"�������QP��r�aH��e��nEDK$"�GQ�����J���A����:`����94v9|-�-���.g�<�'E"i�1W��i�R�\��6�(�s��d!Nj-����
�n�¶���x����+�Bj�ڜ:�hT��K����򭴶E�Y�t�-j
u\S|��B�͋�c:�{�h/�3cch��P~L󣱀i��G��vx����ˢ�$]��1�^�)-j+�鸍�����9���-��$ˍy��n��f<�b���f����u?}���E�Ryh�����N�g],��x�k��+^r�\�di]�&V�� _�#����y��?�œ��w}���a��n�6���*�Á9��{8�%��[^�g=mo�w����(yX��.nhBy(g{=ҥ`�-�3_�_�֍�H� O�~��ي�))�̣"ϲ�5N�`���eh�	�R�m�X�j�<��+2��4:
��
F�K�6�&i)]X����0�	��S�H�����(�Y܍;���:�+Qr�Dt1,Qw���^�^(�N�4Ŝ�3 �?k\����O�ǹ�;&Y���<[��r�����n��~]����+Ai��et��c�}����9���,�4���Cxv2�&���q�~��r'޶�I����ݫ� K�u���SR����Ѻ-�	J�@GQ�]f��A D�eI�=Ǥ���<��Ng&I�R���:���I�;~�$cG��L�LʲIw���(��x�( �E����t(��'ۂ낆�}tW���c+��!��� ��/��?s% ������xh���~�o]�sl[�	g�b]�c+�j��,�30yD��(�x�)�Q>J�#�b��r�1k2�����`��@�����Ű�*-�p^����>� ��������!�X�I��Au����1�vLj�a�O0R���7$]��z�R��d�8�?eW}ƙ�]�f,�p������g)�i��0}h���|�ܵ��0�/�F�[����t�^{��
f�Ull�p�'ᵗ���,�V�®p�_o�����w�K�vs8��T�pn3�b�9��1��#�(�Y�	�߱H΂=;�3e�$��S��9Q�	L�S�c:n�1�s��f'�S�`R���JZ����qZB�͙V�]+��Z��cZl֑��1-ۼVsܷ�
?�vY`:hq<�@�Q�6drIgaRy-�x)���Ĕ,؃&)RU�j�>���ط�ƻ��
���C1�h��m-[�L�'�{?�|�W�Vu�IG⭯�����f�T����0�عk��*e��ng4+9{�8v��8��-8���8_������_?�;���~7~��v)��b���5e��Rņ.w�V1�2�]�Rm�x�[����r13���'�O��~��|��ng��N,5�x��ᒗ���O=�sE_�Y���+��`{�ꖇp�[���Ǯ�1*t���2��-CU2U_=:�4ġCm�\,'&J�t�P���`��j�՚�EĤ������0=�xҺ0y^��Ot󼣧��a#� ��g�@��(� ݫ����8jBM�=��7���9unI/*��|���2p�����$3Iu.tL���rV�h�Օ5�W[6���zϋ�KwV�~"�sa���g����t;-�1s|E�M��b����eԒZ�-U@
7fO�J�N���W�Ae"��Qቆ^Ǟ�䓪�W@-qXG�ѳ��]Z��o�W�#�H�����3ߤca�w�p��YwE���Q-��u�8~��^O�%Z�@`�]Y�h�N�ST�s�1�h��f�F�&=�U	"�����V��I$�����J	���TTeQ��ݖ�t������*I
�L�L2��F�������ixx�p������>�h�΅���M@��]��=9 �g+'>vy��Q�vO������m�f5�&9�~��ݻ�Ĵ��=���/��_|��X*�� ����Z ĠC��y6�l_��'x T�D1&3��tpyG�?�"G�.�qnn�������YشH�B�I;0��4��!��_��gC�� ���O�o��a�iIV��Z�*.Z�:1qe{8ʺ4*�������E���J]aN�Fe�v�3 ^�ӭ� A�cb:�4��n�#�ss��s�[�?�a"��f�Eٕ�3�)s��)����s*̏�G�$vd�2��Q�H���훯�.�?뗴�.۱KqWv�����l�q���Ȅc�:��h�|��2N?�`��w/�3N،�J��ɫ����(����K|��?�#���M+荋�2��*[��c�\�l�3�d��>��	���z���G�7�|�s*�K�aɔ4�lH�6�����(Ȩ�I6��7T~:$s��t�o����S70��:�"鷋�gȥ�#ֹ%��Q f�h3K&�g�R��?vVvbe�c�����g���_z�=t#�Q�P4�*�9��.��knz����]�U6bVjHwZ�r������*�L�c�˽��r�h�ŧ83�f����[k��$g��7���9F�GO����O"0�f�Kd�n�#�b�bXd�l��9C콸.����)�$��m���Y�;�N�) M��T��7�����d�L�5���>�8j�����s���9j[�<����q������P��� B�����Sb�g��>F�ULk�̺8��}p�y��O;Ks�'�;b�v7>�������X�L����	�NG��=�3LA��sR$Mr�(>Z�1��B^�۵
���ʗl�	����V�cZd��~��҈�~LxVט/��Ƣ��|1�����P�u�ٹ,�LL'�c�h�PߚwY�Sy	LG=N6��T���84�Zkar���`Ū��� S�=T&�8��Ż��
��!꘦���'�옾�c_��~�dN9����/U�4���[���\�n~ �^��@�@g���1���tN{�18��`�������G^����;���������ͷ=��w��/ϣP�Xp>^���y�W���[��������8笣~������C��E�h������^KE4K]��������hN���D�'*��`���-��7��o�5}�KR4�u�+QOt^���
�*��()dt���9�ry�2x����z%��"{i�#�h"^9՛�Z��&�GKiR��@�O�Lw�ή� ց� ;۽�g�\EƠV���.oЗ��̙�f^��"�~��ΧE:�3l《e{�2�j<`"� = ��T��n����2v���H�`X7��CvL�[ذ�7�t;m�S��.�;A�|�[�짲V�Sa	V�eM*��Y���ȎFHxq�C���4������K��WP�Ҡh]m���P�m@ c�b�c6q��߁jt.�<�􊮞G&����TC��1�VLc�0�,%=�҉�	�h��ꪀ)O�r��rcf%���
����M�V>2�#Е������ _�o�ʎ)^��ΰ��,-�WT�N0^�"�c��4'�g���tqۏ*%�|�,�n��C��x	N�RV����K�f|�IL 4SpR+����Ώ��ӟ�V[��5�+�疗�a�ݎ�j}��;_��;N��2�c=��g�;�#�!��ڝV��뾭�淯ǯڡ���p�Qy��(i���_�,8%#,��8���q�)��#�~�m��\��uH�M�;��t�F/�C��W�����X�h����o݄���q��\��b�b�a|Yq&A�Q����4���.DR�X�f{Z��bTE�J���#0A�<UO����j	|�3��TO=SW�=��Z$�����*ήs�(6Z 0��%��6�h��ye�A�b�bi
��T�q
�A���.�?(����$��)w�62�;�;�!ZR,�ȓ���Ld�q$���}`a��^Egm��N,�8����K�����.� �3�����	h��^õ7ގ�~x+��F��25B�� r���h�(��Z6��Q��~�p�,����|X�u�n�ڝ��6�Þk9(E/�������4�ד"gm���Ψ`=�A����>Q��������2�7�i�&�0Z+����)o��
�J��;l_��g���u6͹���U����iN�7+��[w����&�x`7F�E�j�/-�{��NŞ����Y�ޤ��U�e�����=�w%�H�R*#��Af�R�-�ZO���+B�E	�d0��o�1~#�U��d�A�faKk7)s[����
8��	L�X�n���C/�)�����S!����:q>�TdS��i^�������V�S�?G~(�����a�����.l��Ǭ�T� �F��/�l��ѷs(��C��:t���0`�|G�?�����0?��x�[� n��C�Z�\�Z�[���N�Ʒ�[�,���{\�߃(
�r?R��@�aJ��kE
3��t�D�-'��a&#E�2.Q�_�`T'ì�B��*yS��H�^A�TƬ�E{�np4�:��4��z�b^�R����i��8��vWSJ(���:';δ�Q���".5���3SiL'}�C���w��<���;0��f3&����^-*/;�o�K�Qy�c���}|�W�݅V˩ ���mx�)G㍯��xڑ؋���3����4x��*�i0y|�+�3�v���!f�9glW�������x�+(Lְ��=��x\L�$��o⾇W�ϗ�i�b�ߍ}6U�in��]�l\���c�BE]��t��}�Ov��\q�f+�Z�UA�P��9�-�&:o&"�#8�:��B������ZL,�x��I\w�y�jYT�����	�Ug�X�J�F3@�����Sn��׌B$8��(�EU����'�����Fz}:�hHUp�]t����J
�,�.8�~�YSZe:�����{1aw�@��Fi��P��*���V����9�V��E4�����;����:-�o����ca M��[�;�%��fؔ��P�x�E�yRB�n�*lIw�:��&I�oЈ�j��*��	�� ���&Y���U%��u)WSIxT����U<RS��M�9�E�b�1W���B}<E��;��ʎ隀i�6�r�!�#vL9WK�̰��Yj�!��k�uD��!j�i~�������Uw�LeO.^L�1`�� >G�y���4��fH���E��x�3�����dNzy�T��GC�QŦ��ʄ<��^t:]�p��h�>M�G�=��~O옢��,S�^g��Ob�z{7���Mx���r`�j������������a�ܵ���k������j;ww�}W�|�\I�Y:���۪�4?b�`g�n���su�`��k�<p�S�u�8��cQ�^��)g��cy?�ů�s��B�i'�����O &0��݀/~�&g��Zy?p�������ݬp�Jn�ħ�+��XЩ���x#Y�\>_oI�kG���(�8�U��w��(%��8�Ʋ$��x�b!-W��VhJ��H�iGȻ>�e�c"�����g$��b�������O6��D@�;��\��=�h��:�۫k�� �F�0��N�C��epg�Ic� E�    IDATh��^Ƙc�^v�x�K��-��D�9���%�����9�K\}�����;��0
6s�ZC��7kZ9�&���v}���!I� ���v��g����lA(޸���._�����ENc�ؚ����ڈ�~L�\�"9��������YAI.�*��b����:�G>g���߁��.��f(l���z�q��*f�6��6�p�YOť>G�Ј+m���u©;��5|���O�z��&E�YRs�q"�}�a�:��.����4i~����O=ݗ��g�(�_��|��L�P{�A�r71x������4��~6bV���2���9�{0iN�s!JB�E���7mh���j���.�b��sϢ|�zQ����?�u41���SLШU�ʕ�
�S1�0Ol`23��N��If�ƑjL)ء�:@�.�l�~�g�A� -@ҿ+���*��jr��s���>%�k5�G.nw$g�I�"�	BH��ɸ��؞WH һJ���&P��H*/g����4�9�0-�9o��9��w��1�q�����������'>����:����;�r�z�fC�tLv�slN�2b� SvL�4c�D�\���j �z�vL�p��`E��-�)eA���q����W���#
w�ϳ7��B`J�fiL?�e|�LO;�昞.`:��'��|���vtZ#��љr�!���F�u�4�!�;@�ꁲ�8��	n��~|�_��;�݆|e�(�욖KetWW0��0Y������?��g�rǩ1��q�ㇾ�{\FnV����h��C�o�U���_x&ڿ)W8��-v�F�3��5 W޲���5x��:ݜ�)7F�n�6����=pĺDD����fn���k�((��� �K39ȃ��5�l�!+����&AQ�I
�A�t�ⰳ�/\(-� }B�1Y����ٍt^�!P*�)Lj�]kǮ�%'9��ʜ�Tո
�cd��������uS�&���)�=�#�H�(�`���\Ѭc�n���fM�H��A��a�byv�	������Թ������lnT����b�:kɢ]�梜�+�e�R;@-1N֋'��UQs�n6َ��:��D&�iƺ
|��u���]Ԩty�M*�v`���VX���]Z���N�~S{�X��A�Of4Boe��Uf<�(7�(4�ҘN�츆Q�#��Lc��W�1;Z�PRy+4?����ץ�V0ݞ�CiLg�|^V}����g��U��΃Sgi�6��?��̮��^w�*��� I A�0"����*b���C��_�߶
��
(��N�<ʨ�@���02��;����pΩ�v��<S����s�w�{��ڨT��}G�|�}�Ng�&Ǩd�u��o�+�����)��ɯ�Ū���=v��N�d�'�/��Ux�2�m��l��$��ס^Z��-\����qGh����m·��\��rO�\��?�u�7�Vk0�5:�;9QE��B/�jkRd��7	3�D�T�|�lFdA�|Z���mX���I����~��8`�}��\9�2��q���o��^���>�>��39�]����q�m+��cyd��Ñ Z��'�	뮕�˨h�1vM��;���A�g&q�4�{jj�E]֡Y�o$)Rڌ��e6��z�&u��h�vLD�� S�����Iw�SO:�)4`�]�+K��sHH�b�+��1�T�6�mZXSŋ���x9�$�c�����IxuP�83�����`�S����Hb+��gq&��ӓ���kr�H��p>}�{1�� ��c��6����㯭o��ۗc���b��F;�S�8�o24T�:Rs�#��"g�U���}ε����%�R�����W��68�]�dE�]'9<��y����?�jRoI%w0@�N��B_8��"��
̭��X[� K��K`���}�����Y`���%d4`�Ϭ%EJ|[B4��k���U���Y����ÑK棘&��}�z!�wJ���Ԛ2���x�����@7U�3IF�`�¶�y����ۮ@:��-=3�����|�K!TUU�:���������alP��ـ
�&���7���{b$��(K���,Eֈ�U���՜C���C�CX�tY�������9P�t�����x�;����Jq�o�h!%�Je�MN�B��E.W@&�qb);��r�BI��D�:������ګ�M{0��1e����Bt%R����^�!f�ސ��������<��z���YOq67�߻�:1eL]�+r\������1�u����#,��,T�@�o:�f3��w�c֒�Sx��G����2J[GĐ���T6oRތ8�v��jەbM��+cڭT�,q�lWf�s�SV��id�(M�|Eu���Z�VR�%�i��o�|��3p�^������������h�t�݅1����^�P�v+�]�$���P����q�9�߿H�]���+*�nk߮Z���9^x��a\�����K#��2���V���	�K#Ha3�ڸ��/ሃv� ���ޥ�Ol�w/�/�4�v�#�i5��l|�[�Ǿ{M�hu�@��F�ٔY����)�ud���G+�wq�ҕ��#�b�H�X�fFjO��>����G��Q��<�Kg����>��$�*�_�4��$�H�y=����X�*�R�YdL�e�����scQB�`آ��P
����N�dtr��wy��I��&%]�#���S��i�Q�7Pc�4?c*�t.�T.�L��*���8��p�k�%��E����f�!NVG�x��9��׵�I
7z_��ҙ��:��4c�s4�I�8c��$��o΀��X�3�t4���#b0��e`ʻ%#Sd����h�GP�9�@��i��+���0`��щ��xUԫxƚZ����xN�U�� C��$�5�k���ǔ�1es?�&�T�9#�ek��%=��jc�h��BF�J�4ٗP�K1h�F��^L̏Z��053��@�!�c�b��uC����:�cJƕ���1�T�'{��E����L=)���Y�@�6�������a:]j[��}c3_�޹��e�β6JmJV���/�����,,�y;�cm �������s���������P/Obdd=����.��g�S���2�14�MT�u���Vk1r�L�&	G�CZ{��R%�JR��0K��t
9zIB	�NTq߲eXv�}x��������,���9�n��I���b�r·߃��_��8M���	l�������G��4��}����#A��.�jc�XZ�������,�\�㧚��s��>�~:98�^+M����8(�y�㖩��3����@�3O�M�)�~���d�1�$1��Ύ��h�Q�+<\$�Jܹ�Y��%k݌�4�+����9!��g�G�ܽ�UϾ���d��͂;�Cp_�+A���K����:v���Y���x f�1�X����dј����Ϭ��7-ţϾ�R+�tn@<+��8Rj�LYM�C6�Z�-T�x�фS �;�����p�>����ĥ�˄�դW�Z�\sVY��ԃ@VY�� XV\��g��!�J䬵9��6��_5�	1ϵ����,�Ocw���%�f�4e=�lS=-��I6��S3��6&~�:���f�VY�{]�z�ab����$r�\�����e/m .�����5��h[���sbB�ڬ�Q����=Ķa#���O�S�"+\���(h��/Zï+���E�P����]"n�R��G���F��s�����Rib�P��V�g�<R[������lUD�T���S�ܾ���}�TKJ��i!�k!��"�hJ���[�j�6c~�tA���7��"A�	�����6k�6����|���7�"1ԛ$v�HgU�Ù���|N~ɔ<7K����)6�@߃�
%�\��`̋r/��!Ҵ�,
*k�!�B)�4JyR|e�$1�*zZ��.�,��[*奪O&c���d�eg.dӪN��֜I
��T)��؛Re�櫳ݲ+悔������a��aμ��i|�JMT��O����4���T��+����������cR�tk{n��?����L[�^�ƚ�w.�#�p���.�ow����͕��G1��f�\y=��)�Zm�g��O>�<�$̙�w)�e胃��S+=��,f��!s�ï���V���� ��8Z����Ibs�����Ñϗ�%�G zb��F�yeD� ��8R�&����[��^��ke���қX��Q��v*U�Y
�f�ı���̓��hx��~y�#X��҉�V�|%tK��,�ʼDޱ��#�j��Jcx�k�Ԁ�W�%`El�E�ʍlrV-��fR��r�q�LZX:�1i���KX�P"ͪ���E�����T�@�%�h2�Tg�90U9FZ�O6�R�J��8�����rȊ�	��q��{��W*hQ[O�bѼ'�$���"��ʞ�N�x+?V܈�����+�tV���Uy]T2s��duT���++72{˄�6�*=���9�y�W��Z���#R!��y��W�}t��V�]��ww��J3s��j�2�Y�'���"=8��lU�j��"��'�R��n3.)b���/�X.���k�="05P�^q�~�!s��l.��L��"V�Lu�-��\��@\��4�h��K߃�f��3����3A%c*}�d�#s�b�R��%t�UIp5q�dƔjՏwAM��p����&Kl[����w
v�G��F��.���00��{A��������ǧ�8sg���0�<�y��o�[F��|6�zu�[ףUڀ;���?���%`L#�A�9����T�"�J#���j2|zQ�X�`�Q���s��ofW��>�����^��",�?��b(g�ʛۖ>�?/}JX鏞|_�+�	&�2)�&���~��o��T29���9�I�m�2.9��QS�H�$������N?&%a��6f���h��S�a��یi����)�g�����&3v�"�-�{j,�e�HF&�0��QArԯ�J7�����e��|���F2� 	��!��;����ac���1�^ٲZ})���+>��)����*0oF���8�]{a[��M�3c���j���q��˰��Q�@�倉$�ҼH<��Nց�(t �qS�K�дo��SʜL�b��l�ϓ�k��0�q^���}�<#�o�ZUwu���J��SU4�'��30�c�nz��zPh��n���a����=��uk ��p'Ģ�-����;��m[q�"3�f�*q�Q�i���⸣��Y��}�B���e$�1)�����ϸ��ը��n����2��\'PsB@%��ꆾƾqh���ËLQpxM�������a�1��b,t���׌��zP88�� ����cL��˔����0x�~gJ�ھ=�q&Xa��� S��]����}�nX��t�����aO<�
ּ6�D��#����:�e��ޟĂy��i� 
)�p������I�}f�K+����q���0^[?�R�4<�H�B�����	^d�A�T��C�)fV�䀳�~/\'�c�4�b! ��3-_��!0MF�i���6�PTh�9��0�=S�C9�$��d�@�Z�Ô�6��0).ۮ�V����BB�H�Dsx���2ZSg�gL'4'��GU�K�T��l74e��0o&*Q`� �UdZ��{nZ��Kv��ld\L��e���z��m�����֥�%R8h�����%����W���_��˟�������G�ηm���c�I{�ա�AN��LV9��+ƀ���������Q���j��iN"��`ִ.>�<~ЮV�Wk�܂���f�yyX�?�G����a�>�pɷ����I^¡���p�wɏ��-j�nˠ�B����߃t�0x��&~�X��8���R�!��^j�Uv��$�}�X$c��c��DDjhGc Ұ�EL�\�k�����!7U��JR \1�G_1��bN�k6��xn5Z��a|�"�\��H��R��0rfVu�4`j.���2Y�&r�D\�ʓe�\��{�R��¨��+��V�)3��_�Z�����l��S2gM�n% ��&"z��`�s��)��!�Fq��e�&+�[ AO*-ϰ��k���L�)�
Dy�-�����Ԩ�C���ؘH�`�H�0rH�|.�|�o0����Ɋ��E�Xb�G ;�l�(8Z/�}�!�gg)$K�1!��0a�s�g�Am�T
ٟ!2;5��"M�So�>:�v���m39��y��1e��2��
�s�s�~W͏8nF�9�cCfZ2C�e�c
�]˄@]y��J�6߿#��W�!��'r/��}I? ����V�z���4�O}�hs��(&�L�+r7�`���t����J��U|��P�$Qm�0ш�{_�o�x*�
��(�L�G6�Sވy�]|�����beJ�`/B�U�T�e�Μ���~�e�$>�O�[���N�V��>��jB�I�Iʕ�z�i��n�-4��]���|׃/⦻����#q�~;!/�]���I�_ޏ?��Z���E�
Eq^�\=e:�?/�)3E�Whmo�ȑ ۖk b1M�S&}D�s��:��	���l�)��1]+�>m��:N�p�L�#z���ף�M�+x���/�c��9�R_ρJ0�Rሂ��P�E�@��m�Ar&�\N���j�$�*������T�=]�����G=7ܣ�#�
�v��(f;��N��K�W�y�e^� R1&�����U�܅�66�N��g��T����7~V3<]��W��j�7��R>��(�1�2��^�)��a��v�d���S�F��zYm���W�Βgc�d�CS-�Jk���
Ly��=e
�)��-j��9ik��]c����w&�5�O�I&�?-X����V:��6k��M#�+c��w�٧���@�8s$�:ë!L;�2b��~q�]�����'���)=��t�O�L��ױ�!<�ȌBɽ0X�,ku-���L�=�QK~��|��`3}ͅ��a-O�Ք"q�u+��F��T�J%�4y���sn'�{q����.w�����u"�_aۂ�D>����b��5��u�i�c�݆��/���g�$A0Zx|n��qlibd����[U�հp�A|�G���ܙ1q��:�G��oێۄ�����\w��c��(�)�-"F�0�6a��[�%��y&�tgP���a�,�.@407���C����C[���j�Jd�{[�^�NWSq�%0e�3�E�d
]^�K�(�V��L�24?J�����0̲��Q��ǔ�1��b���f?m��!��	��
Z�Z��^g2!>��W�9��$�*kx&�=c�,랄N�*��|w�����;��������ǔ���\}�}2�����P`����?���^�ŗ�˖=*��/~�c����T̈́,��@����?Za�֋���7��
~�۰y(W����ՑIV1g0�K.8�-�5Y� E)�E�]��/mE�����d3m,�w'�迿��v.ʁ��|���῾y�X�mS6��z�V����m���c�,�1�z���^�����ӆ�H�D���Z��O�.�9���JO�-�(��c@��{����XSo���8��E�'&^Q��f:�B��C����n�]7�FN�ıvxdc� 
�o�/q���h�%Jb~D�;����G/�F[*����J�J�4��	c�*&�Ǽ?"�m�1m�^���5A)���� 6����k	��$���RcԈ����ofR�1�,
���r��dY�?L�&��|):?`Y"�5)�(͑L�F���JuHXrM���0���S�����z��p��UE��C�C�S"X`��80�V<]h艃�&-���Әb���5�%��Ћ�R��t=��g�@�f�4��+ ���4U`�{�����R�λUk�16�&���T1�tN�RSr��	J~ɘ�+�$��%	��[CU��>d9.&��̾��;-�x�L�� �최d%�&R^g����\.�y	�z�(S��2\���7�mw    IDATgR@�>�=v*�g�C�E�(,�r)�H���|�xq�z̝3�E�i�oSX�������
����l�g����0�u:�M�eF�?��8�����&�4���^}O?�K:s�n$TΙ��
��߶8�u��;���Pi��ųϮ���HzK�N��Ҡ�p�`�e�x��Rq��)G����s,���8\���ko��t��
V\ݐf7YbL�#3G��J���n�p�q!,��=�LS��O*�;T�VS؞�}(EC���wϐB�p��߰w��B>�K�L���oի� �e��L;�KB,���=����+�=�������SE�%�X��T�Z�Z��� ��K�T��"��:f/ou������ ��})�T�W$�Иp��/O�O�?���k�gf�M-�	�Y��⋠�A��9#�ݤ ����q�i��L�\N��P�U-�}��# ������a� �O5��v�k�L��,��P2�Z�
�SȨ�Qv�8ՈE֝ʵ0��/?�t=������5Yc,pˈ��wAT��,��5,�)��h�a��t8�!p��$:��2��>�x���E$�#�TGz��1��F���� �xp6��e���f,P��<'�sV��:���/�6��@{tOzU�i3#3��޷)���h=�]y!��ڼ�f���h�UK��A6���8���2�j��mQ��u����x��Z�
���U��-��F@Es-��WP|�Z�:��y�&i�D���;lO|�Ga(��|�)��n~}�c��_���xUL*�h`�@g�t>t�Q��]i��F0~���� �z.�*P������yw.{Õ8��Bi,��2�j�������4����
��(�W�90U,�렢��*��#�I��3M_�'R�s�R=��3בִ��:锌�!k	�H�ccL	L9ǴS�brt��5\�R�<���~U��*�Y�$�27fk�D�JU
���k��fd4 ����q�8H�o��\6F�-Pbtխ!���;��_�(�ٹ�?0��^O��2��o�_*���>���݇dp�\���*,�Q�����|G��/ U0]�V6�*���Q�3���Rފg^iಟހG�\�J� ��^��l���Ӂ��u_<_@�$� ||� S2���[�˶q�~;�>�=v헞TVjּ��\{3�]��*g���e��q�9ga�yC⨵����:��O`�hži�f�Ȥ('H	(�������n�L�Y��%$l\ڡ`�z��ܟ�&p�G������w_�l6�Mrѵ�M��L� �J��V�h��I9��׎�b�үX����NrDW��t�w#��D�$�vX6ZM��eT*e9����}}(�E�+���4�֛���S�g��ԊfQ�I��H���V��L�G\�oX�Φ�?s�$�%��zC� �XB@�Ȋ��O���*��&a&�ʖR��}�j"4���G��Ii����Sc�)_�������=� Y�AX7��i��I�B��dˌ]�H�����]yhI�L�hA��������2�{%��Xi�>6�v�!��2C����@> �,x(0�&z2�):�rH� �2z-��H"K`:KS����%Z�膙B�����$�np|�LP��s�I3I��[{��I��N�sB���"�}�{�_�:{�:��Y��`��cx|�j�ݴ�,~'�sg ��c�o�w<�Ǟ\�
2~��Lʆ��G���b���/���*�,@k��|�zx�����3��#���PXذ5��,7D�&2��m�TF-�MLl��`��f�>�־�'�|2r��(\|v'��'����"c��Y'���E�I�J
c:\��{q�+�NN��8��)C�	�
��4��Q��R�gWQ�~2`�E,�]-�8�M⧲����-�c"%��@$R�m�oS�A�SVU�DљSa��PcId���Ti�ESi?~��P�
��|�ͶAFB���3$��-��D궱JS���w�s�*GBѡ]�\�x1���Cus���}�=x�Q��!�}��q�51 �����o��Z�4&��{9�2�XJ�(�� �4�����sW�(��_�4�:�d{���s�#e2�����$[�CXx;w%0P*O�	����5).�$��&�m���@Vh��E%e�uKh�d���j�pyJ"�j*��4N!\��������p,�78���-	,�SX�f|e��Z��-4�0=��g�>'�;�����ts�5��M%�7����<�r��N�i��f"�����(~f�y0�S*4��Y��!ܡգ��23
�g��e�M�!0�`�}?j���s��Ύ�~�\@��^�K�9RH����׌���66����|�ׂ�	sW1"jw�����L�c��W>q�2Z�%@c��v����w�݋F��n��'���G��3��.s���Ӵ��O2�ZZ�����ݙ�I�2�XOb'&E��6���a�x��%�M��I���nU� �)�}�ʰE=˾�&�I1��τ�3��ēC����h)b~��"<͏zb�)֧�d/��Lh���j�$-f�'��^c����hQS��l�>d`�,�>̒����Le�=Jp-���)A�Ǭ����D� ^��ҞѨ!�q1�,�?���q�c�LG����V*��m>�=��s>��ΔEAM�S�m��.�%V<�{�:���X�c�̼s;�����ȵU[�#�'�򾅁暇�?އr-)IQ�:�|�)�����3`�W"K�����\'��'Xir�B����칠O�y39K�JU�^A]_��\�I�~�WJ��\���|[';(��P(��(�cC�ѐ�E�+�6aN�e� dE}=�,p��*PF���z	*�A���XBM�q1p��^?�*�A�ɯ�%V����e`��Q�se�44�H6��HPБL�h�x.~!Uj��$[ʛ�Q-�������<�h�֚�O*�K�"Y��f�b�@ds%��C>��Ι0�"�Ϡop n�N�r%���r�����W��?�]�:�ɪ�Vq`*�@ݔ^��>WM2�2."��B�I�\#I\R=%�E�q�7�4�M�wB�_7�>K�=a�5)k�oOP���y:d`t8�ϊ�eRH���f�(�:/vեY^��E��a��EZ�����L�2��dp��لZbq�e�K��	t*t	L�)d��#=��LRX�1�A$2]@敁6FSaL��wOH��l_ɟl��\�fCZx`�19���7d���~'��ĩ�;�(.��-`��������`�P��?�9��6��{%�y�T�$�}�$ȦS"�V&0�e=��^����\�
�Ɍ˺xq���n\���k%���y"o5���k���P�W˒p���'��94F��/�Ö/�.[�S?x��D�&_j�(�k�˸��'D���)/e;Q�����T�tN�:2�T�&�>��"�#��b���m9`U
�)��Vޞ�s�����F�E$���}�?�FzW�w������Y6�O)8PV�9�ݙW���^M�#'��]8`5��4��)>��A�m`6��B��ʀ�+#g��I�}>�o�)F�G�9Sf�s)�*�k���)�����%+��G��߳�
�Ȫ(М֩��l�7��5w��1�H��`_!�o8t�L���~�:���xaH���~dg�M��l�R��EM�k��G�P�CI[�A��*ս�앢�������fN�cM��3�6�Qa9B��g��(u�gk��و"D�
>��{bh���1�sj5������e�j�bd��2�)��6yۨZ��\ݫQ�Z?�4��L�-g3I�f��n��zy�NO����Y��.�43�4�rP�U��s�k�~7��^�8���t\M�}�}>SUJ�!�U��<��pޛh��D���a/,x|p%��_`����𜷞hgL��Pp�2S�(Ό�<'���-
�9t�Z�8�Yϫ�M��@���3�)���yg-���o�4-}}���Kqݭ��7I8h�y�ʹ���)��Sw��B���gd99�%���Wtb�����a)n��S���P��70h�?,�GB6�=F��8��A�.��M����$�%	F�@����D֫��1��k�<��S�Vkcڭ5TMr� �3�����k�r}2�W���n7��&GFd�:��y�g��H{L��!����s��#0������1c��F��2[����s9!.�tK��Q�6ڵ*�q1���t����a��3�X����z�ȭ5��K�`���p䒷�s��'�`�TC脶b�:\|ٯ��Ï��%{����G����4�3�c���ni]��낒�t��وo�jli�4YA�]Ɣ���b�1�a5���6�K��q1�n֐�u�ǂ!|�3���}w�Ț��L���g��n�xx`M��~)Y�j�������ʬ�N��VKei�Ɖlb�j,A�-zn��?�*ޑ~l6�M���gUd��)�q��Y�3_����0ȤZ�7���nz".nr������5�i^���M�9w��\V��9��Ԩk/��O��l6����ep2MY�^u��Ҋ�ZG����hqI�
�`�d(l��TR��T�@n"5� ����V��l_}���ֲbGF{rx\d	
J�0����D%3dL�5%qԜ�$3�3SE�Cb�w$�Z�O3R���nDD�0�^���a�J��jt�h��|��ޝ�Q�V�b`���H}#_��Y��0�>�
� �Y��lZ6ԋ���(���#0�G�4��lV�%��i�������IzC;=���ɘ��.ӕ����0��H�k�)�[��*'��/^%��F[{Lk���lr*R�!�jAzڤ�I3EQ��:��m�ئW�ێ}��i���w/�@��V�<�?ݶ<�Zƫ��qƩ���sҘ���~9�����}H��'�W�\6���F��h#v���.�
��;W$���ѓ?@
Zm<��3����D��${f̚�Y�'�����>���$q�QQ�Z���L!E7ӄ������m�x�A�s��8���q�QG!N��*m�1������'��q��8d���U󣘸�^��;q�]���D,�/���S1~�#��so�� �5�gf	����GY��og&z󢪁 �z�T��E�`k��p��T]w�U��Hd�v�O�<oE0����^g"b5�`��6�eaJ��3���8�*;�΢��&�fV�uoI��n�����]zB��wL&n�ۯ�c�3*��}o��F��[c��{�çN_��
*��dY��0�^\[�U�܋�X�R�z�~Ē47"��@B�(Z���!���@�Ӂ�[�����w^�5�2#a˅�����%��
����A�2hk ��6�5�u��lj��fB��Z���|u��p�K��`ᘅe���i���4ө6�E��.ٚ��#d���X�I���G�M�i4�b���� ����)�8��}A�6�ۇ`N���A`+\�$e"�mTP�؈��GN>
�~��$A��n{��E�� ����5��mO`��wV&�L~$�
@u@-V��3Z��QG�M��6��Cg�=�sDۼ�١��5v�{<	U��*�7�B�qEU/Qc%:@��ȃ�(1�#E4��H�~ZT�=#���Ս7u]��M�vu$�t��$0��ؽ:�	�uҡ8��`�>D��$��v���ޅ�n_&g݁�\��|�=8d��Qd��'���֧)V�c���,��uW���_��O��e�r�d�T*��0)���e���L��A�IݰM� J1�XV`J�d�0�,��S��L���,��(��D�͏X��~6`�I�e�i�k���O2 �JƔ�G}�4�2rK�������y��ɡE(��e���l����� �v]"���I�*�&b.k���b�1M*Xe�Ml�Zmt�1mcz�3��m��?�m��4��/���m�ӽ�.2`���So��˯��O<��O8
����㞷Eh�H��75o��{���5�[!���������"II@|�͈�{(c�z?oO� r�|�G7`�+�2o��i �l#��b�=����Y�#�s�rԂJwd?�t3G�	<�r	��a9�>�2�]�*��L�=��˞IGL��=48׳V�%RR~@�0vmu��c��r��ɍ�e�0�Ҫ�v0I��/�Fɖ�0f3Hd�(���(�-<�K��2������ZtΗ��F����ԼV�T5���"��+2X=���N�ʘ(M�Z�"�N`��Π�9+}3�?�RI�0
J�\ds���Y��T�DF> 
�
�ɢ4(�t���|�͜&��F8#㨌��1�TC���ʌ5�%�$OUL���/"27G>ў�Ps�ζޖ �5�Sh��M�cNgr�x���im/���լ�kg�������Ҵʥ������$C^�5�szmLO<!�����a:�D_�t̈́�^w`)�3n��M4h`$�G0��o��^Q���NYJ�9����U8Q���5���&�rn�db)5�hvĕ������`E�B�3H�ͳ%�H����:���Ϝ�w���x��~+��nX��ZC�y��O����� w`�kM���`�����P��_��C�G�0mNn��9I��.�w����I -��W<�B�a��t��Wwe�+��S���0��������II�,Ϥ�E/�e�"C+W<��_��v��#��.gL�Js�>qT ܿ�M���G��p扇��vDNb�X$`����ށ��~��L��d� �i��2�Ajf��1}�e!rP�K�͚�g���F d#E
�$h�^�=��q�M�X�1U�g��Ո�����|�d^ei��5�Us5=S� Q���\ng]�g�9�2|����x�&_��QO�=�֘�Lh��)�
�8L�]$��fa�_?�!��N�/}{nIVT�'#2րλO<?��^unZ���Y��$��S吶���J)���b��K�*��;�"G>�H=�~k�&	�M��[�^:�[�$���g�Z�퇌(���%���(�{M��@��B"�Ԯ�r�ao5�5x2�7��^����ޡʁew�N�z*)��T���YN����z��QD�㉑�ru-�L�	%��C�γ�}�{qԝ�u�i���V����~Y����xӪ�Ѫ��SA.^��8�=�d̛d�(I�`+cϼ\p�mX����6��C͜dd]J�2���~�z��v|�l#V��[��C2!�I�Ц��e��/T�8����q�P�����Ԁ�S�i-���-\뽏�\��S������6e��3bL)y��[/��Zﴐ�֐l��'�Ϝ�?S@�$���_�������ݹ��o���Y��+3�VQU�k׏��u��h�Q�TPoT1sƀ�
�e�,ɨ!+>��D(��k��2.�������TSHԗ>fؚQ�������n��2�3�GZ��D�����
L�;,N�8��mL+���fh���'3�q,_6�v�`�`[[d�D�<{HkU���Ь�Ӄ�$'R�d^{L�ɧ1��&��eҒw	�P��KS
��\V�Si�A�ܨI� �h`�F��1mI�i��D����9$�t�ى�Y�K$O��[�����R�,�>xo�����A�"��?�W��j<��S8�����~D�x�J�C������̶c�5&p\�ol����b�So�:�D2�A*^���wϟ
LYY��(.��MX��0r����'�m���Ʈ�p̑�p���E1˱&m��5��5l��f͞)���Ưm�⇿�	˞�F: ųH��b���f%�#����0�
�&i�C��JT��Vp�� ��G��"1L�Ó(�ڰ�]+��>'�ȳg���D���#�bpD9���	�y�)��X���⿩�.�z�-��h��3�IS�ʃX����L�&i9�x]�F'��hՑ-d18c:�d|M���^��+���kӹ��d�z�Ȥ��f��_+�tfb��ބ�    IDAT�����"���.
���fsa�&F�Q��T���ȩ3oF{g]6fR^Q���Iܑ��{ES4k%_jp|+h��K�S���(n���
�u�\h4&�*�v�.5�)c��N�&�w�⪂Xs�uT�Ł�+A�Uh�+x���Һ�Pf��$�TGG�F'���43P�Q1q��Df�8����{l�rE�5kgL����`�Qp,�YT:Ɗ���zՆT���27eZ�z^���˒L�u�n��5�쎋����~?����ӥB���>ܳl%���]�W?�O8r�,��̃rxx����i<��z��i]�N%P���u˛�T6c��� ���N��c1K�_�U����0m� �]��X����������V)�P����T���TJr�
I�sL%��1M�FO>�(��.�0o'|茏 ;Ч�/q�"�]��M\w�ra��>�]8t��5GM� 3@̿����v�|����I����zK���;��A!���?j�/hq���f�&����3�a<�����z�]0��G_h4v~�����y�%��0F�8�Lj���L*Q3�*PQh�u�gd1E*�)��ɭ�/�B�� v�wtF?_p���n?b$��%�4��y-6���(�:������6�o|�8��J�'J�W:��m�忼	Ͽ6*3+9$��ȱ���H�&��vt���7�Զ��fx��N�j7 k1#(np��y��:k�ʎz�J	�Ҥ �D���B.�D&C��/z��_�����54}�,
������\#�>8S���:h3��b�1�ce��W0>^��Z��r��j���r�.�lFf�Dq��p,��"�͋��.E�:?{O���%g0���eY"~�ya,�s++"2�W�n-�xR��S�����V��Z�-����c��<��ir+����"�X�zߺ�v<���n��<K͉��O��nd�L!Q�e�� �>�n	-�E��&�^>(.G������=���l%1,����0WS��? ��E�PmgǶ� ���U�V�S&s�v�D$�=C�v�n��>z�a��i
L�V����7ʸ��p�+�x߽�9���_�
ڕ��Oڋ�o��?�?��0^xq�����k�7���x����N<�>r1��)��B�<�c1Q~>�J����xd�$
ӑ�ăE�Z���ն-ϋ4�
=:�y�(�(0u��?���B�BQ��)�T�@LГ�8�q1"�m�S��X=RiKJ�{L��4�����R��KC��b:���^CISz�t�HfC`�Ti�������
�H%0�+����td6��4��	oe-mmq��KUէ#���H�Q��L{G�5$�bv������< �ԁo_�\w�r�3}����Y'b����x�>�ʁ��8�C��y�|:�oI����F5Ft��6��ۿ˂v`�8�����G֠<^C2�E&QƜ1\t>���Wt^��������r������	�8'��޹3N8�ݨU�x��W�r�j�R	���c��-@6�m�
��ww�ƥ��y2�V'�}P�0q����$9��3��������Bͦ��j���;�<�+&��nY��HJ��t6UK�j&�*I8�F���}}�6�R���ã2'��I�h97T�l�֙�5L"�I+�/ +%��՚���ɸ S:��/D��na|bR�)D������!��W�q��d�OC#��I�E ΊM�������	��A�^���$��K2�V*�"[Rwa�'JL;��E� c���19>��(�iKf��1��	�)If��I�{1�o��Jrا��痲��:z���G�+�Se����~���4����SY�"3���y>�������y�ܥE��$���f�w_ ��V��\ ��=�A�>#��d�����]^+x��OɌ5�KQEz� F��6��h�k�0����`����{���8��DI*�vtM&0�M�C����cJ`JcV𴗚2�8gb!IW^Jd��z��2�Pޓ����VJ��h�I�L�VB�Y�P_������v '��?9�������y�i��;f�p���{�"2I�m���[_�nX�n,/��i�UÖ-4Vڈ�����[_���	�< ��2n��F1=:��å`�ɞW�5�=��r�.�*���h��V�d�B�Ĥ`���q���c�����y��I�o�4���^���,����r�{q�>;��!3�qo��pѕ��֥���t�yq��b|�8g�R.�uG�O)^؛zQH���hH8]�Fהn��E���;v�B)�D����1_��,&w.�p��AO^�9J�"�$M��e&8��z�}��L�4�F����uń'�!�5��;D�}�%"̊���]7��qg�FkZ�I[/��);�R�c��I|��g`�l�\���Łzx��-��;��K[Q���M�w�U��RgJ�,c��0���7+?i,�~n3[c�｛�pit���I�r/I���[m��5�j�&�ѮW��wj,��Q,���;vǂ�c���N�+ �M�/�E_!�~���7�1n��K��X��N2($�T�ZR���r����
�xs+�}�u<��+xs�8��V�3EĒY$�.�e�$X�EiM�0E��\��Y7���!s��9�?/I����3˜x;�
:M�DlE1Qŉ�,�g?~�M�"y��-���ϯy�{�%�yrOx��2-(�G���9�����8��t[���-q��}7�-� ��e�Elf5��}�9�A�C3/�E���B�D�)�q��6�?`���U��x���'��������~O��T>C2�-�
2��:)
L�ͺ�^����_㉧_���s?~*�{�f@�/��g_؀���f,}h%��$ZȢ�H�*�ZC�]C*����"�;� |c����w�'`�$��{���7�އ^D"?فA1���i��*)7u����e�K^�d��U��&Y.�+/�)�_�����q�ٷ��R��q1�&MGC`J).b�Ⱥ�'Y���3���Q����4#=���Ίx�*��oK����N�c�m���!�ϋ$�����:���p�*(5����F�V`���Ƚg�睅�g%�w"TcGcZ�=�ցp5��s��&�dO|��`��3�a����g���?�#�y�i|��G�?��I�90E
�	�6��$V�~[��XL��h��?�>�&F�(dH�&1ۀ�K
0� c�Гø�7���JD�t[������q����|4�ʣXL�Tn�λ����pN>���'!��
Z農����n�z�@r:��ˌL2��_�65"I��T��C���T��֫&����»�Iq���!�/�?�U,/�F�����}��@MN��h�����'�^t��x��s?19��oVzb'��Y/WP+UP��������J
0����Ą�a�M��O0MgӘ&li?���Hw�cb?-6���H�'F?����B>���A����2K��Pk�02:��[FP��L�Py����ЎuP��/=�)��tژ�@ilR�YIJ���1M	s$ ;-����Wdh9҆F:���ٲ%LDN!�S3@�D���U8]n燸@�#������+�AUN�	����:W=���O�'��d�;S�:� 0,�5xH���������2�4��1`�e4?����~�I��jS\u�e��8�%�� �Αq`��G�H2�I&�&��et*tw�T�-ޏ̬~t2	aW(OiK0o׸�V�f�J�ZS^CX(qcN�9%I,�{jO���(��0��(l��w��,�c׼X��֭y��������*L�:�(�c�5#�߷�~��nfF�9Y����	���: 5�[(�nTD��(m��Yq\vѿ�w���"��^q�>��r)��h��Ͱ�14�Ф����~���0Q�-n�z(�l�x��q�5�b�%8����.�Ș�u��x7����>}�q8h�푑$��B�xs������yC�TV�R*P����h��ɓ�9M"d���0�e�Ps���P�o�����G�>���J<Z�a��8���8g�^s�f/Q�4�[�{8��Qp�qY��+�f~ �h��{���P~���ЗX����͡X~��a����Iw�$`6��o�	��Ez��>�.RT��'9]��T��Upʱ�p�c� ]Ӂ�	������K��z&'����3���f�a�^�X`�L^a��'�xf��j$�5^�?��2
�TQ���E��@`n4>�FiM���#��Kb��|eh�{� ��?� ̙�d��9��S*J\e��"�@�Àx���v�	�D@��&0Q6lncœ/`�x�ŵ�l��c�C�͛dr�+\����ZܐujRl��	�%���P��`��j�5_��˹e�_��f�z�����:Z�	����O���;��O��w�%�l�X�V��;|/mh���&�{�o;�)��҃J?R��k�˲�bg�����/{h�z
G�1�aÀŁ@��k6:�V__�jj>��}+d���rT�n�_�yq�s4���wǁ)��θ?��n���y�V��y���Č�������?����]�gV�����}*�9pW�g�;�����׷��_݄�r}�wD�o�TZ�����qt[U��%MK�+��(�8�HL�\�p�W6���kqߊ��K �?C�A�+���}n*-f�M��W�Eүn�達�v\��5� ����3���5S
���mA���T`���Ӥ��!cJ`��u`*�PJ5?*�)�鸘0��I�YԼJx�gL�m4$W��� G��Yek#�T�9G�iޤ
G�`ڒ�	�*�1��<�,,R)��kQ��z�t�����Z\�rG�6|�c'	c�UY����ʵ��O��?�w�N\����t:�M1F�~_�����0u��(y�%?�	�>��R�^�dC�b��/��%��͙�p�%��6�n@�V�T�/��/�ˉ8��]�����s���[������n�:��8�5�_�ep�o���76�+�i���M�O�􊠆��[Փ1eO%YS�#�5u�j�T������L��g��g�yXŔj��>qI�����0s�$�0������O�)���"8z;���;��'ШօU��+�{J�VCȼ�ӑ�l1%|�|���1���i��L�qDL2�z��C�h�2��C�lC��x�d�\30�P���a"���(U��@�Z�R�&��l@�����´"R�A
L+�e�3�=�E`J92�y�&����iwѨ��꽔�ٳ����i��|]�wi/�IB���)k����g��˄Y|pv<���0��3b�a���pk�ӓU�D˜NM(����)�N2��\kE.�BD��v"�X1#�)T>#S��Q�!���i��@k��f�&���L!7�����t�ӄDg�	�P�x2��,��e)jHa%�D~��t �L\̘Z�7���PH3?g��1e��H�}��Hx��а@��>&̺�9�]�o���Q�܈��6��?�NV�g���a���/�6�r��&m̜Q@�=�w����s0o��l�j���-����#�B�˱H	4�%�o�t�=\��~{�C`�T�L��`��P�����<AP؇��J~�����ɘ@�J���>�������G�3l͕�O������k��mw=��p�G߇C� ��)�׷tp����W��Q/Y�FbI�g��Պo��)2PgJ1�a���Fr]5�Y�^����B����R�L+���LP`���`Us-8�M5�ۿ[b���k��gL����I�'Ķ�l̏��pg��5���:ɵ]��$�A�k�
�p|L�&h�w�RE{;ޯEc4����q�1{��5'1�?�;��@_��݀��܌v,$������";e��~R;?h�����2J�Ay��U�@Ȓ�+*ͶbCpo�5u\��t�γn4Q��@�L��Z�q�1��B����#= ��;����@��8�����'J(��v#Ɛ���>�8`�Q=I\�jE��C�FU���5�-���GVឥ+��ak�f
�L?b���"r�>�AN%�GeHTƭ_V>q�T�[(Q���4*�pU�TE�J�ɦ��[Kzy�Y�dɡө��(!�e�Q�V���M��z���R�^��L���N7hU&�� ���zʟ��|N��$S�?!h��ב���wT�e���ճ��Tu���{$���R��'���vض��'�����y<^	�9o`gc����l�����%)C�7�e�>�`���0��!%6xIQb�\����㩕kp����O��w4߀)WB��կ��-[��r��Ll��B��Q�Q�A �q�˨�m@1��'>r<��/��i7C�+�V�m��9��&坁��,t��Č#�u' ���}V�2��\�r���)�����-0�$���c��L2�|�[�8����I�1���e��.U�Θ&RvM�+ �g���q`��)0ͥl'G����}�dL�Ƙ��Z�T��\^='r9�5�NUj�#mN�1��&d�0��2��N��'���6Eʋv��8�z�,�c�`f�3��^�Gm>��]~���!W�������g��<�Z7��W���?�}�Q�s��Օ�b� Y6��j��
L5I��o�|�U��*p粗p�u�a�˛Q����6�&f ���y8�`��z�e�3c��������j�
R��3���O����Hnk�����n��z�	��g.�R�4p��$��=��Z'�T.���23VL
h�D�&�NG�6S�nr�JBl�rx�_���`* P���[��̀�W�]*T0��f��T��	��&��Vk�R��ā	�#�k:zf�9��f�j�ݹ��C��##�q&%�;$�Jc�7b����C`ZC��B�����'=-�u�a�4��g�h8�%~V���(}�"/��]&7�d��A��>��Y�%0��4�G	Pz�u�Y6��Ia��z	L9΀r�&3A���e=��%l�Sm^.��f���5��q)��M�(�f��,�In#;ĥ�^����ʾ��l���A	4�{��E�I�c*{V+̼m�����"��:��H���OΏe���J�	&�c�9ns�"�)��~�	��V��o�T��ZQ`ZGslR�)�E��b��0��Yh�G5�9��g*:�]�x-2r�%R`����c�Y�dB- Kna��SW(?K�G�UC��K������0���u.�oVp���g�_�J��gmN/��.���×�=sg������w�5h��ыg��K���@���W~�?�g`�K�Ҋ[w(�t`*IN<��̙eoPRg��`EZ��ђ1]Rl�{b���ּ����9sf�ͦ8�)�tW���^�4��p�iGc�>�M��n���?�}�U�c�*H��x�	�ʗܕ�
7j������d�٩W� {u���A�踿M��ro�M��"gde�r4��}޳�'?�-����3AZ;匓�4�_�¡������Z2Z���&Mj���������	T���/�;]���q�<����j���s^gݯ����9Ec=L&�6����2��-�^	:x�8�q�ϒEU[�N����9�j�^d���!�"�vvT��,o��c�@n)<�zK����s�6��%�r�Յ�*Y��:�I$:�8ԏ=v����/~��<��r�� rG�U�s��)s~���\�U�����ϓ���|�);�L^��A�ً�,��������[��ɗ�����k�Q��Њe���!S��L�fS
Py��`l ԕ�V��1Aһ��&�M�PVAb��lo����=�2֦m>���4�$��*�FMF���&A��thz��RC+�������G�嬁qSpN�QW�k�V��L�h� ؑR��m�����l3yA9\�d}]8cJݻ\<�D�~ۓ�oۘx9c���гB�=�6S�ip��=�^����K:���i�UF�W���/�>z8�]�1e����X��V��~�ǟ|G��=�C8d�9�'X@�Իl��v��    IDAT-���Q��2�5�gm/��j��b� �c�ڗ�e���vp�����<	��H��eX�i��x�:�훿���mA,;�3g�]R���聢쯰�qW)(U���1�3��1�)��K̓L�6ƋEQ�5�n&�xs�e�<G6�@�g�S���	EBpʶ9z�8��XO1��V#���e3��t�ݾ��E�XD<�IJ�K�Vy�W`�E���~��Xk0�#A�%���͠P�^�y�n�L͏�f�e�%z�8z����������M�;?�7������n8��c��C�5����X�y���Ë�����	Itt�h]�T��O.'����Ah�S��5�Z��uŃ+^���	�������÷��\y��b��}G)��M��_�U/lB�����0��]�.�Ƨ�pG��2�t�������ӎ��Ϟ#���cU<���m��1{�(��p���U7>�r+�� S�W��0���� �!XsY(?'�z1Kx� 49y�;�hb��
0��������oJ*]=G��$p1�vv�������6:t�e�W"���Ae>O팺���2n�Vb
�2��H*cʟ+����l>�3��1���y�O
0�_��eV��8�F�S�)ʱ9��F��*���L� q$HPP�C�=<lɘv]�
(��3������DE���W�@((�s����O�� C�Em4ɘ���Sc�
���M=�S�)�]R�ʨ��8�!;Ēna�WMGʜjFeǑ;��%N֑�z�	�{���q���'��Ɠ ���I'����l��U+r��㮫
Y$�
HO�C'͞S�G��-�m��O��=���K`��G�?/���wut���$�4@ �(����|��2� ;��Sm%�ت+�$�ƾ21"0Mp*�i�.=���S�$�����Y�:a�����&�nVѬc�������b"Qs�&����xs��t1�S��l�0g�t��\�}�9i���GK���kQ��d('�Bs��׊�ю�m��үa�=g(c��P�3&1Rm�B�L_��$�#�m��gVc���eL3�r�,��톆���zh%Ճu�`���m�|ds
T5�?EW̉.p�����e��N�qƉ�`�;���Uk����6��፸����NH� N����G�7-<-�Y0P�
��,�ig��AVh=�7N�n.=r��������5et�F�Uv��m�]�[��9v0���zdm��3�!H2Y6�9gC��3�(��4�Ԣ��y�P,�Oސ1ݶ�Q�aO�� ����,i3��A��r��H��c��2��+�#�.َ�S��\�6�	�6�[��XI7|*#�q�x+�5+ף9	�7Y}�ʃ�C�s7��r�ByՉa4+���J�&�X��,Y��u�"�:�{��c������8)(v��/Q��M�;�M���,kۣr\�7�v�6
Z#��=	�)��$��� ^z��O����de�5�*�[7t4MCӤ&��("�~"��E�'�8
D�Q��GPPT��349�����*��Y;�sn��=�O{��{�N����k���~7�� �{�9��1$�s�.�E*?�#g�#���;H�gM+r�H4s��u�+@�P�Wd^�3��>�a��Ŗ5�İ9�,��W�'�ݐ�'$SH��mB���>%"B,�i���{�d��T3�o�O���_�B3�����#���L�M����S*���3����yA�Wg���fL������C��+l���?d6r�$��i�1P��q��a�tЭ"�+����~�1���R�"�ǳ/�q��?ŝ�<��9���i8p�)��b!�����	/nnaޒݑ��v��z�!S&�:2�y6��,��e��'��,�Ħw�W��:�������� �E~d�8W�D ɗL�(�N���=8D�e���$�����xc�4QT�#�P���b��2)đF\&��@�\A�*���+�c�� ���W�7,�K�TC�4
����&'�n6e�%�id�
Hr$9s^���I�g-�e��dL�M�I���� ��K�)���r�l�����$�I��v�(`ǭY�/~�t�b���U��P,`Jg�+��G�����Yg����+����|~��R�}�J���O}g��x������G���ݦ~X�ں:�e�l�/��:�����2����◎�1g���~�c8���f?�`v�%|��WⱧ6��`zf�C��G�o~�؁�L[=��W������>r���\w�ݸ��?ǧ���:d������O/��A�,��$(W�@l�%�f�$H3i�~S�:�h1�n�VW���AJboö}n���f�d�S�w9��$D��f��}���5	L���H���XI�(+Б>=��%�a�����z��
j�)�L��� S��)W*
L�maS�Ο/=��ߴį�Td��A�DN�1cjy�yVd��xH�	L�h�:r��1v���6Ac]�cp`�C,Gn8�\�ݴ��d	��SU�,rne��a�˚�/;�!m�[�	��)��W;�,�屬�J�KW�y� ��B�?jI�z�H.���̜�����+�@E��J��Q1��i	��i�M�Y�i���Č`_]�;-V��g\S#����0k����0#E�����r-��� ��tx�9���KyHK�+�7RDJ�)����HzSD:J�V\���@��Gt��:2��s�����&Պ�X�j\�Ύ}��J`�*��9rf�<�-��GB�Vkc2ה�.%�)8��	���N©��a�Z��&��b�m���������'��ע/�KJ{@�:����4Ʊd��}��ww��Ez�ej�&���rIl�2��}���Km宻b�8�Z�.	%�9���f���F�{19�FG��n7e�S*��ః��.;/A1���@��ӨV�߲UzV��Ɠ�xɈz�D@{L	Lo��9\s�}�$x�;���{/B��9�6w���[|��zd��
����j�5�����w���b ����o�ˀ�t�e\�(���Κ!��~>�Q��e�r	��Ƿ���!0����'����PX�z��5�*��e��Raxr�)��.Yֳ�I�uIr��
�3��=�Z��7�[o�{�é8��f�ӫ�L��~��V��33z��r1���ؼN�~��w���:��\-��Ff��X"�����sL�E��g���G�>%�}v_�c���'vY>�9dG�H�1���[�&r.��f?��Y�����up$ͳ���W�S�nS��;Sk�ʒv�~*'j-`�<�nW��6<����<�B��D*?��B)&e���~e�#3kÖf}s{&�nL���ђ�����\�d����DBi3�e�����g����WW�y��_����}_Hg>r->�Ӂ�][�D��v?���+}����V(R��?�Dy>Ƽ�k�Qpv?����Fu?��=�h!J���|�>0�s�/q)v��j�%�o��2p*g�
��ܫ�i">��������<�c�<Hլ�P�9��7�z/;� ��'����,@�m�����7�q��n�շ<�nb��9�R�h7��4�Nb|�z�lz	K��3ވ���h�+�do�<d �<WƧ�p	�mj#���LaD</��@dc:=CS�C^@`גּ�r/�ҭ�̎��,z
0�"
Ly����������ŭ� S��N`J��*��Y��>O��JΤ��L ��O'e�)]}Kʘ2%M��-!A9��8h���
�T�R�R��A����j,���sL�i).3���K�%�z�lL�i���H�r�i���b����b�\5?� �΀<���Iyyۏ8`>���a���	o �g_�ƅ���v��&��c����!,e	�XS��Z��&Na=� k���
�T�����<��������.q���B*��h���~�c8��=d���hV����w��x����xMOoCa8���������c�G�#��̳�c͞��Ǟ+�����n��|���ƾ��He�f?��Z\�Q��D�B�:JZ4ت�W]�4���mRgf2���izJ��m�I�,���h獏"0	�-|aX-Pj�Qh�6�$F�U�᮰�T֩?��6ָl��T@�_�J�8�q+�1ԪU���E�N�S��|��Ky{(��Ny��j96g挍
k�i4P����'�xDaL�Y��)!R<�P��C��ҊZ6F"�\6+�nx�)�%�+�*�妲B��p�<g�r�m�05鰚��� �Љ�Ys9	�j�ZS]	]�a���gU3�+��μ����y�Vb=5�V�����J��ie�O��a��=�}���=�Xɋ���d�JU(5��)�.����<�v�%U6V��=��b���,��c1Tk-t�It�i�Fǐ���Ȱآ�����^��f�(n��� Ӧ\C<��Q#�bKnX��QHʖ�]w)/͏:���zD����s�ŕ��#�ɐ1�`�� s�R�>�,N��[���k��L��Q9��9�(�C(c��f�x�n�����55�@�hE�j��/�B�wl�O}��8�!/O�8�Ri��1hl�c������Us@1���D���L[�NJ���,�-�݁��} �%y��9L)���z4��TmI��Y�r�rt���>��Ʋ���s3��W����2m�X�{�8��ñ`�0L+�=����_�u7?(܏���S.�>��^��~��^?�2ފ9�w���s���$P�㻪F,L�R����
� x���?�hK6<�S���CXb�=g�� ;d�n�s�����*�!�RZ�#�X��|+_��g ��S5�(aX�k�Sw0�}e�8�{��h���Duf���������R���ɯ.Z~;��<��s7'9��� B~: W&Q�d[R�=��K��tཱི;���U_�Lv_�W���Z���&�
��$p�^�q���}v��E)Q�s��M[!�9׬�GO�Ur��D�P�s?6���Vm:����~�Y|u��Y��K�$��4�g�\�8���8,��Vp�gɽ	
�)(�5b���ֈ�*���&���A�z�x���Ty�G�AJ�v����p�?}�>:ͽf=PF���W��**����,��;�̚!�V�O[���=/��Z��5%��`�/+dY��oЪ�#-H{�	I��(W2��F��fY�A1YsB��f;��3[�Q��Ȭd�;T�����`�����gcj�ϋ�h��E+���+X�
H���앤��N9j/|��o�|����6�2���_�n��A�����ރ��7�IȾ���#���}|
?���X��6�� ����t&�F����Кق5��>z*N>zw�.��@�^>5��|��xu�ʎ!�.�\t����έ�4�t�RA|^�33���/ʘ�!d�=څ�敢�fc~$�4&��&��;h��I�7�W� !FW^�Z�����$Ϡ�B&%R^���&'%���g!)���r[Q�Q���^3�I��A�4?"8�xJ��B^��TZl��J�)�u`*�"��cʼ�����.�`�wvb���m-������N���<hw���2\5���K�����;D�4��+������8�5Ȉ
�dAa��2�B	[������������K���4��bF����1�i��'��X��9 z����<�����J�b8��]��s>��L���՛��,�FG��^<��Q|�cɈ��ϯx�^u?J�pL
�n�1�����Ϥ=�ҿH�ʤ��pʯ�����к8FE�W���Ī�R���퉎��2��10R'P)SX8�P������ٟ5<:*sQ	�+�2*3�j���i� ��)YU��J��j�.�)?���(�F��6ku�g�hSF�Q�sJ�z[9��+�7Ai����2V@�3e:��)�"�e5FLn�?���lR�t�c}��&隨����IR�g���F��3���1T�4~j(��A5�&����H��� �IgDG{I��w.pX֊�&�v}ƌDA�}4��\\�kɀ!���dQ�l����Sb@@������g�`�j�*Y�:V�X�]W,��yE�!3	��M�X�eO��Ku`t!��6{RY5���}雐�|n~u��zK��=#E$������=9U։l�Hy�+�7�\Z�L���`ڤ4�0�2^s�;�q1t�%cZo(0��=�j�dg�Dq��[��-v���}�YŠSƼ� �zÑx����96�;P=����:@h�g��K����$FP*J��R�2���M�7�b�9}|�[�ÚUc�n)�׊�'��W^-��R�<R�&�Kx����꘮�РiABg��FK�Q��0Q�ىPe��?_�- �b�6�阸��2�w�&ݦ�[\��z�~�s�]e$�p1/�e�(S��5w⾵O��n�#g�	�\�%/l���߹w>��Ԉ�1eEV�zb��%�J�$�qQ���#�<hϗ�;9P=��%ճ��א�g�H@hQ�؟Y��&�	��H�L9���2#�@,�W�C�u�V���{-�j茣�H���F �,fĿ�>wx��F�=�~�D׬���Yާ�`Co�����_ή�����C�9K��^�s�Q@ʈY��<bU$y"�3Z��k	b��,���*U2�T����B[d��P]�!�����z�V�AC��k9^{ľ8d�]�tA9������͆�FHB���"��h`�l�:�M���W7㕍[01Y�b�)UB-��w�}����x����,�(�9�-G*���Q� �Q��X0o�7X�+�����qKL3�2�4�j>�EF^3j�	��J7�����Q<��ڱ!7C'�T��iR}�"(��ӜkMJ�ن�|j��N����p���e�r]Gtߚ+��G|\���
����>x�H��^ŸW|[����������y�v*�ߞa��ŦY�MH����J ?�B׾)F|�:h�k�ס��o wP�1����m^� ��}68f3F���Q_I!��*)�GƔ=���$�;h|��NÒ!2��:�8z|�t�Op�=��>����w���F
?�=g�[K�}+~u�b�7:�^���S�ЮN�]ڄ#��_������#�#ތ�h�t����^��3��B?��G����u��v�q)�Ha��,깥m-Ѝ1���]yY<�!Yn�gq�{W�)����k���t�դ���)A.͏4N2�(0"0���Rީ)�ϧ=��b�\FS��*(��3g3id8���C}rZ\y���HD0e_/q�Ǌ�LE���I`ڮ�߮�]`����������ё��].����v����8@��H��%|��Wছ�A�4��B
�~ۉ8�#������/��&w`l�Y�f��ӓ�B��?�_]~&f�5H�����f���t�s^G`jۤ&����/�
O>�M\e+�i$���R|��?�����NP�sm��Z�.�>�F����C&�{f�ޯn��w>�z'�L6'	{9�Y�����.��W�q�f癩��Fmӭ�t}C������\O9���en�J5�(!*y��h5O�B&c�Y�t)�j�z�|�fP@Y.OpS�8L�t����IEl(}�I2�Ğ ����A�T&��#Ø3gD�Aa�\P�}/�@q�(��j�I)�\M�w��Rj0'a������Tm:g���J����%2I�4�⽷9�USiX������7�ZeȘr���J����t�| 	�H�<k��fP����U&Z#�!�ϯ�d�!���>*�Sl9{�H���P3#,9�#���Na�M�ѫb�hG�揍�Պ㶻��ƭU��:�Y1���q<�ZU�z����؁:���q˃O��uӨ��P���M���^�+��4��	�I`ڤ��ɢ�O��h�aV ���y�A(�q1LK�t���F�F���[���+e�Li������Juz�����5Ȥ��(��k�i�F3�r)�)2TE��9����M�C���9�g1\P��H]]T�vJ��m �x݃���(W���02\T�>>@�Z�����V�`��9�s�    IDAT���ǚU�b����p��a����ӣ!����#��c�_i�"��![��f7���J��t�LfO�_�N�����4~�y˕=��f�V�M��`�\6���b��e(�2�x����_�j���}
/��"��i�<	��\�_%Y*�=�ۿ�]�n� ;�N,��4����7��K���3
L��@�j��R^�=�b���\YA��F9)��Q@�";7����9�:Y�a�c�_����Y̍X�V}浨	Z�{1,4!r�I�,�EG�yg`�?�����TŤJ54������#2fBf���Z���Π�� a����h�`cD�J��X4W�Q՘(Dzh@Y�=���6�D��h���썊K�ŉ�����j�z��4b�i�z1N}�18��}�x.$�%�s(��W�-A\�`������2�Ͼ8��׽�M['�����2>�Z��z��F��.?��{��Q�,��3�V~^&��^��n�D9�� 3@̿L�{Ȧb2�f���lV��'v�q1��dJ�T<8��\��&�Ң@��@��3/U��?ޅko}�*@27�d���ేMe�#(l�IAix%M�kz��A��Q<�E\ߋ���6�O�����?-��hO.Po�FH���^��"���%�N_}�(���-��WI��s�ҮO��l��3 �?ώo��}�ά"�v�T=t����nT�Y��mMi��� ̇¶"1�ӴL��DxK-��ۭ:��
z�i��2|�gb������-��O�����v�ZQJ�d�ϩ'��9sG�0������I|��ߣ�-bt�21G���D�:�Ԡ��D���0|�7`٢,�� ��������y��jg�~�b��T�"��p��a�Ձi���c� �0*đIy�24�6�,�XN�fw�
L�M�j5t-q��5mR^1Q�RSz��/��]I��z#��dQ����I!�H��	L���ʡO�|L�~a�\��i���I�LӅ��2�{K���R]�#�{3?�{d�����kR��5q�٧R��0=�������)R���+>z�[q���֌��nK��ᕸ��031-s?����g�z��4�9lgWoB	��m���>�#�� ~������qV9��|6�A��|�&����� S�������߽
Ϯ�����Z�v;--����S�;;-�k��ޖ��ź~��Ǟ|�V�]vB�,t���:��˿�ٗJhv���U�+�Bf?�={Z��*��ژ���Gʸ�+�4k��ʹ/�}��9�H	��D�6���b	@Q/��h� xkr`������R!2� i���>P`J��tJ�E%��6(��k�g^g��1eՅ#,�i�F�F0glD�ϕ:��l6��Z"B�#a�ؓkUV���̗S�E%���C��L�.�����!�� �� ���Q_����_��JbĞJ�,�ySI��g,qT�@�R�k���fb��<����2p~E�
�n������~0S#Mb� �]c�m���fL5i���"�#,���W���M��>���f��(�M?��><��˨5[X�b!>�Σp�޹��k��Ɋ9��O��۞l�Ow=��_-�N�U���Rq�e�� �j�+��������dL�_��{��5V����r��
��H3 ��f�0����)g�bi�!!@4�bGՁiO��(��h����+��hHϒ-]����-4[딑���t�0V�K�Cq� ���Kݷ�y�6�W����[	�!��I���d.+�i�lیX{
��p���kvV�����ڜ��㡇�@�RG������B�T��j`Vow1>]ý?��n}�.g4�d�ߟ#"Ɏ
;�C�=��.ұv_���v^�P�Jb/N��U�?���7�hwz��02\��yy)l�	�J��������=�y|3���F/�x:���	D�b��aQN7��
L)��c �u0�2N��U%N+�Y�u��=�������˓`��WY��q�՝�2O���p�&�*'�xnf.�@p��ΔYIQP�R�5/��j�Ec�,̀%0�	�뀙��9D$��b�cN�(KA�95Q0��/?g�B�TRAo�K�Qj!�U��Q������,��'�/�vWwܮ Wm�Q HPJt[�5�h��`�Po8� ������
��ǜ�h�s��I-�U����>y�e�v�Cx���,�ʊ^�m��y�$VRm�e��E]���g���v��Щ쯮;���y^j�����6�.�:�2:�
��.�-���Q��Gv -(��$�g��N�t==ׯ��UZ�=���ˮ��k�C��E~t�����l3�S�ْ��퉿\��Ko���DW����iG�/�~+�k&
F�W�ם�/lm��E:\0�^p��� 7P��Gg�����Tw;�s�QA~������~	C�����ul�[���s��3ѾV}_�[���+k�k�A����)�մF���v�f	�NI&||������h�Nxy�8.������dl��#^�_>�_�b�yHĹrh�����8��o\���~H��7H��y��*V��;�p8�x�츀�� ������ݱ�_����h��_J��g�^���@�a�ܿǿz��+{���W��-hT(+��T�z(c�P`�h�_��S��I�,�ǲْ�J���2/������4����<S��JIe�.J�)A�������P�N&��aj����$���`��?0ƴ�>���	�n����ʌ�&�'T`u�iU�%,ߟ�s?y�ߌ�	Q��ۀ1�9���-�p���sw�~+�����Z ���$^�R��?�
7ݲӓ%�x�bM�^��~��8h�J�P�M��g1�
�tIk(/���n�p�/�����C�N���ؠ� �edU|휳p�	!0e�|��������KH�SL[�2�6�]�������#2�.��觞�ĵ�ދ�ׯ�k�?�9hodR@�\u�+���`��
6���f&s2��27y���;�T����X���C)}lrv��_E}���)�V��A��v�.=�E�n&M<��L�V��J��d�̄�GȘ�N'Qo6Q)ql��VbJЗ�2���Q�6�l��l���udt�����ۑ��V���-֙d3(�Q�SȤL�,��fGϑ5A������i�EZͶ�me� �BV�Ǵ�W)o��D?L�d�z%�hbL��<hj�W-�P-өTM�h��nX��*������/L�J�9�[3к�n~OH<I�����Uh�w-�.ꇝ b;�!�R���GG��Nc��+�t���ꊣ�*�.�7���<�S�t,�|��o��Ok�FY��7c1��~s���˽���ϣ�J�9ӕ�L���ZL���d��"�&�~	���* -�&z�Q��T�"P���E�1M%�ǴE@�ĉfXd���W�8g�V���BL@���1����X��>>7Q�u��O��,H��^�F�
��HrPn�-���$x�!@"���/��!�+Jؠt�!�����Z�F�4�doK�z��~{�((c*{F�I���p39������k�*�e2���?W����:�B?�S�?)�i��kI�,eoq���m|�C���߰�)�udA(�D�1�FT�t���E���Ε�뱍���ѣ� e�Lf�I��_�'Z&z��o	��Ur� IWȉg-&�t9h1W��dv9�yt�8F���	�V���Z����'�z�62ÒIa?��	b��l���S��ǎ0�t����6�+�o�b}��g�?D�&r�-)	h��Y��KW��T���T�l?���v��������Jb�l�$�Rp5�rݞ���|��Ք�v�4JېT�z�(�z�x��X��$z�+�THf�2�Lg���L���p�=���^��T����9���A�b��ͮqA�l��x�eI~�Ę)Xd�\���F:���~��������k,�N��,al$��[�#_�?=p/�jƆXP��+�еa�����ƭ���=�koyO��D-�BaQZ-x�&R�5:V6�K #kɀ��g�E�$����ȸ�v*��Qx!�O�a����s�y�"���k�tF/ˣ�����]��9m���S�%Q����)i��ړ�5R� r�k�9{�=�s6��C��1[s�0EcV@����w�Tc�ͩ�Q�	�F�a�V��l��*�Ӛˇ��s?����P��Ź��n���tӝ�����+v����%�Fc�&�G)l�P��^��y�e�:�Bu�L����3�u���}����h".�R���nǕ}��4��h�Ȃ�,o�S�9P�����>'�~S}C���7G�DM�'�o�����=Vd\��{'0%[�Q-|��f�Hi�y�2A@so�z�����i�#ku�4\5`��d>k��l�R"���)��z�ML�S�s�{��,��<zT!�׶��1U331��k0��%0m�� 0��w~�?�&�8x�]���B.	ԑ�K�k��Ϯƍ�<�j���~��|����]���|�}�X2?�M˽��@q�P��֐y��Ɣk=l�2�{���(&�]$3E��5jU�8Ⱥ9�L�����q�r�����;��W.�/m�bxh�Z�A�Lé&��/`��vĮ+w��d�s:�}<�ĳX�ؓ�)�`���pЁ�aΜ1T;	�����`�¡ϴHת�SV+tn�U���j��!R�NfD���42Y����FSd���Y��q6,s�.��ϣ1����2��"�!���S���J]�`=L��|k��bpD6��Y-7  �ە�Y�e�W0��0�d/����5`�E��@��2`j����xsf?+��θ�:�Yz#�g��p��1T{r��P) MY.��	L�J�OW��Z�k��g���łT\Ӵ�p�V��R*+��Q��2�ُu���"}.���FH��ꎕ o����9;�ײy������_{�BO%$]���z�*�q|��*��t8�v�=l%�����Q����.���k��3�L�񩏾��?�K�OH$�6Gc�1Ԥ�Ka� ������0��I����<]^	�D�[#cJ���MD���<���V㊔� ��ƚmtKet,��wL��ܨ�����M5�#S^{=�3�`��&b8&��gc��}P�׃U
6V�f�FV0�V�o�c�d<M�rYZ�m��i���Đ�h�4?O.[�y�4)�s	��T�z��8R�2��o|{윗�4b_o,�ƕH>�"�/ǿ�Ui�������2м�B����V����o�q4��[����>s��8���®�x.`��lG9.�����	`�
-���_��ϸ������Z�R����U�Ӏ���k���ml2��~�X����i�������'�?Q���>��Q�/ �NQ����2��l�-�Qb�A4j�U�#ƸF�P�GwgR�4J���V���q	㍎���O��wU��ZLf%���,�sM럡�V���b�g�m;�"�&c�)K��g���e�5 ��|��O��i[����O1��H�K���~<��;ݭNc(��	��ƻ�x4X=v�/�j����!��G��]>�G�|�'k��G@1�4�<Oh� <�8�s�ӽ?emn|E��c���EM��C�>W}Ttpbo�1�"m�u����۔��k�P+O�Rs�|�����#��I��}W�{c�EZ-����β���u=��7����_F��E<�l��T��\�������F���c���*ҋ����l�h��d/��|�u䦂�K�`0�S��lY+�I�<0'������pF�'Q���_����D�Y����ۆd�՗�Xj�4^82"Z&��%���3�����X�u�Z3nT���pj�#/@�c�(�U_�ݗ�/~�.HH���������1�2I���e#f��r�O��z��~����Z��9���G�8+���p�������}<�T_�����8�͗�Q,E�Y{Ȗ�9 ��̫%��������T�]崇␌Y!�*y����MӘ�����2�ԁ)Y����Jq%gO��" �g���ptzbB�A]�K`�8��2Й��O{Ȥ�(c�EmbZ\y	L�`N�ˢϑ5�9�<)8nU�K�W�����dL)�=v�E8��a���B�5]��(:�����[���?�p�������;q�K���7���K���<�F����"�ل,<�d,�a�XkV�SN<
��\�]�B)���lY�~�_���4�V7�J��r��j��X��Dz��2�f�'Q-mC�5�4�8�sƛ_����h^t��p�E����i��倽W�#��	���赫xy������~�64����:t`m�0�Ū�wŎ˗#�A+='[ز��n��GdM�mW3���c׀����>���i6K6/+����Q����Y�t�ҾSI��dGFj�l"�{��+�[h�J�tV�C�or��a`$r2��ȉl�K1m�6T�^4���|!K�ܤ̹lT�Ju8� ��ǜ9s$�k�-�q09mû:��Hnh&G������.�DZ4kl���z�.=��Z}�r�rC�w�K�?ke�,�K��=σ�RMJ4Mʫ��TKU���Z���!!����e<���y�k��wt�v?��Yj2�4�S�V��ڹ�Exb�����} T(8M��vc��G|��ފ9I�UQ����s�>��G	��Oc���g��ҧ�}�7���=ٴ���x�	 �>8�_\�6��\j��6E�T�i�F�R��1�%ui���!�<Ä�����IVޚ�`�)wJy�sF��;�n*.ë��7i�����$YW�!gou�7�#4�[�� R���f�:[�_U���o�I�i|�תTm�<%K�|�:Z4`o4� .=�\�,�PZ�'+Ϟs�n6�x��m�����V��X2��k���W�!k��#cb���C!�+�4���ًI?ط|-n��9tb9����`W��@)\��nm�����G�κ����+��¡Š��M��L��q�?��>�"��1�;4xH��
�7_ح��*
:B��O�D�i&d�/�u9{'r$ڏg�%W�������=������(�XZ������ŮkV�hIs�5��� a7s$3��D���F�y �?�w'ƙ�9�.�@��K��R,�$�n|䝳
�%fy���ܼȍڤp+G��E\zÜИ�H�����������+��~�A�>w)@X���贛h7��4*H��X�0���vN9f/,�tK���b�'nB/���i[���8��c-�yi�v\>)�'i&dry)��a�g%ﳈ�Y03�?�8ғ%c�|�_�x��.GZr����_�������XN9siJ�Z7�Zi�F	�X��p�A{�-�������e�I$)\2�Yn��a𧛟�o�t7֏P�/��H)�F�TR�6����<4i�~���2
�ռ��N����V�ڶN�1�������(X��i�������Bh�k�=�ne��\cP�
�W�~�uE�O�$kv���"1Q���&[�"_�H�^��@q/zG㉉�݌Q�Z�cb����k��rQ���G��¤Sc�����]�Oi�"���6��o ���~\��?b��i�\��������Cn<�����m���>~�q����'�H�-�
\c���3�}�#Y��bsͭEA62F�w�@�M�������4U���
L��������VG�ќŘ��7Qȃ΄���!�2}٣d<��Θ�}�)����
0uW�dRf��)��Q����1�	�tRF��-3��
����� S��ʸ����`��|����b 0=��o�!{� 5�=������j�t���z(�bt�6�7��5*�M��[��Pf�5{�c�8�W��!��b�5Z2�ॗ7Ⱨ���=	$$rh���')u�Q�|Q��d�ʥ)�����do
_�܇�� ���m����|�x���9t���$q���24k    IDAT��g�����41��ߏ{x��g��r�1,\� �q8v�q�#y<����_v�~aZ]I�$�
�z��K�6�<9��4����JJ��^�ݳ��P��ОS�	% ){N���M�l�0r�\�9���$��8��)��Ѡ/A5`(i���W޻C+i��pv(���^+�#3���O�( 8Cn(�|>/�"�kt���Q���l���L����rF�%��f=kn0Ŋj��io�ۖ�%`fo��l.�DZ��8%	r�Ǥ7�ϵ�W�%)%ēR��0�!p��o>��
4s*UU�Kpe�e0gVX�1�L�L�킧����\Ȧ��cb"I�&�"}�D�����z])z�hU���MJdf>�ס%�JE���/j׶b��C�ޗ>�%�)���}��ث���E�:����X:�E��}<����"LNM�g'�t��	�� �{h���Il�� �V4��������#��tF�er���\]cT����A�)sL�ժ��Jf=��y��	cG��b6����̥t�v9.�'�t���V'0c�˼g�m|YC���%~�X�Y}	�Sq)�p-��Z��#ǁ�=�.�@�ss}�n�c���d��(��>U`�q��3��Ѯ�c�(p�g>�C�,�Jl��Z�O&��B��!��G�PY:<��B��}|�����u�"���E2�R b���m�D�1���~=N<z7sr&�򴊫� �6#��:]�!�%:ڳw�<�l��<��6ĳ�h��q)عT9�gj�Iz
��&��mʠFYO����v3QFOo�'|Q�љ�hRU�菆=��gg�<ٓ���m�-?���B�j��|�'�n�!���vk��ju�]=�@MA��`�PU�ʖ*$Aw9�9��}֥ܵ�b�0�Z��ϫ����l��;������W-�}�����o��l�e�xkc	�PȚșh��x�j�Ѫ͠Q�p�����	g��8{�bh�g��FO\�2/���M`��2�[���	<��T�I4��bY�R�YU�K6��T(jϤΘ�K�t��<+���tLճ"�]�읝�~f�޷��dv?	����R;�h�`�uDY�$��fe�T0���7��>k��	ƒ2�O���?��H�ӯ��n�{+~��7���M� ]�{�z�h|=kA#zf�- �(4�i���f����Ƚ(0u��`����������Y����-_t2`{#JQ�zHC���>�������zU�cJ��Vv
�Y�}ܗ.�7�"��*�����7�_ [������c Wb�2��q=K�1�à]��s�����	0����j�糖� x�s��ڔ�����ބ��Gx��8��58�?������[�s������f����?���������C,=�d.��W����,�S͕�X��g�6`Ե@$�9�e2�,�$	L)��k2$ ���r1ޓ�X���{L��s���d���J�Tl 2�(0e~"-a4�V�T�DY��1J�]dS)�Y�;*�e�)��8�
0eۍ�U:0���������r��#�v�~��$��g!���{�j����'c�A������+7��}wQƔ�	���ٍu|�W�f�z_�����B�h�e�P��k%1���1<���pQ�r�ZG���2.���DZ�v��L���"-��d������P/s.�$�)|�3��O9P�d����ʅWʬ�D��7M��&�ڣ�ƿ��d�0Oo��֦m{	�zKg�; ؤ��8ĞB�xq�֏��{ۄj�=Y*�%�JN�T;w����pK��^�^�����j͸uM��i��QLQ�j�TA�S�*^�Vi�5�G{$I0)��`��<��(�p�CO�XM�tZh��RU��S]t�h��bO��FζɶT63bz��'4C.��âYo�C�E?�B�  �H���gbWg&J2�����`���F�0����ǯ�U��d
�7�@z_�4|H���gڢ����(b\o1�Vέ���{��A1t�!_,H%�<S1�#�hB��&B�%�~�١Co L=�����b�S}�z#}��3�Π�9�RQPj���U�1��	�M�A�(�3�O����{��g��a{/FΌ@z�l߂�?#�X�>*�~���p�w$L�?�>���`��`Z2`��??�M�4��Np�AB�)���h�u�)���"5�G�3��-���4_	���S��SJy	<y0���C���������q1�����=��fG@�S��c���W�s����s}�Ñ�W*��g����Lc#�*���'2���$:��1y�PfO�J�-�k��x��5)��!^)���L���Ŋe�0o,����"o��dkN)�К��	�	1�:�@�T�<��K�ˍ�����Hg)��W1�Hj��k����b�V�8��w�'3N�<Ҍ]ң��#ö�~��n��ҁ�q4[1l�2�{�>��Y��� ��9�X5��I&�R��Hĸ�y��~���FAM��cc|���,A�"O4Ե�oݤ�co�����:��Gu�$\M�U���A�Q�*�42;NH|��+�9���o�8q3՟�qR��:����\&u����,#�FcDM�-�m�G��/�O����iQȁ{��
����<����K��0��^)�hҪ"֚B1Y��_w(�~��m�!����O��D�6M�p뽏�ֻ�ϭG��D,SD��,��NI&���M�n���ݝ�%�3F[��߁i '�����ޙ�T�G��7��񳆋"hKg�:�
��j�I���H�j�q�0�y����c����}Jǌ���NB�i ��X;����X��$���q橍�a��˽l^�q~��E����@�������Rt��V��v ���X�?�[	�V�.�`]���E��O�-(��]���m`���бX�`V��E����#tdDJ�ꬰ��b�,�44o��3W%,��L��UI��iaQ��R^�ŗ����|{,K;ȝ�">+(�Z���U^8�ǡϤ9���n`3��?�/��w��X��٧c�R0���r1`�\ۋ��7�ō%�z��d�2��U��b������!"K)h�
A��4$�D�''�8�-KdL��t0�5A�+�\ĐĐ$�S�U͏�	!��^U�9ŀ�M�b�},�f1�D�y���2G�����Xkκ�����)MMSb~D`Z�6�[�T�$����$��BsP�a�Hzk��Jy�BF`�^M��1{/��g����w�ts��E��?�p�,���]�O|�T��b�M$� �kp�m��ӊ�8<���1uR$���N7G)�b���K3^1vH$�1&Dt���M�Fyk����d�Mc��� �Z�A�2�ze��i�����S�x� S�"0��	�w�xf�4:�S�/,����?��,p��\����"c��s�����	��K��M���j'����|R�����0_�ȋ�z�T�]R�K�[�7�#'��������} M9����w')qг���rBa삀c=Uf~$3�x�E�)��RH�k�˚�i2ƍ�j�06��n+wĪ�V ���7p�̺Z�`�ݖc�=Vbт1��U<��&<��:��t(�a��Ģ�sd�(G�LN�13�@.?,r&&�����$��2�����j�&�d�2�v�{�H&zb��ϥ%��ql/�#� �C"1��yC-ʆ���`j��\�Ip
�xqff%�O�������>�LR`Z��W0���nd�h���;'D��G�Y݀����,l�ѵ�I�xb�22� �TO�0{8��rq7Y8�ZA{#�e4יڄB�����P��ԓ�xX�aɻ��1�����}a�r��N=��X�t����cq�\}�&��ڧ���D�ϙ�,&�GZ{#i`o�Q�؞ZC{2�cHs�&L�GS��$���e*�6z��,`J��tq�ycʘʈJy{A��[�f#��Ȩ�~��8g|:0��F���ƕ�fŅ��$�����VX���ּ�=�M,Mc��b���s9L��x�ōx��W11�E"SD���{q����Z�nS���F��t�e$���HJ�\�6i^��TU�"�ӞA"�� Ff4�J��f/��И$�	�5S5�\��D�N�Y��:��:R�
�4r9���ɚ.����>E�ݡ���&/�|�r)b��3�i��d�T��ǝh�n���1�\zRN9�&�����_�Z��1�Q t�lQ�0�(��>0=0l����t���Q5>@FOY�ޜ**<�3�0�Й��>9�tp|�fO>�8葞T���R�(d@���"	��*���&��z,�$?�d��������7.;�2F�O��xt�G��5
#��� ���I�]/!�)a��>�N�)G�t�=i2_[Z
̉���v���ݟo/�c��G�*�d�tN��q��Z>gu�g�Ncw8FL
���k�[���41���~6������p��(��h��#-5/����O��z�X�.2��=���̹2�E��l��U;-���'u ͡d�r�1V�q]�	8}�ɺ�����+�ګ��{~H"<\Y�C�,����L�"�=&Rm�I��{������^Q,��F�R^��c�X�`�Y��
2�=hC�f�,>ȧ���@�)L�ֲ��"E�����`�����,��Y*� 5�sW���S|a��3i(9�GS�Il�-r���������!���i^;�����E�C��!�'�i���u8�����m�8���ދ�vR`*�'4�n	���x���H�&Q5�}\���M(�K5��;_2�-�*��e.�
�s���)g�J�m����X�&0ͱ���U��K9����5*�b�,by�C�1բ��[�0-OO�`��c�i���f��*3�Q��/mE:�0�V9ϊ���)�E�K�P5p
gn˙o��qD�IzZ����?���� SNk�A��g�3�8�=��_x)�|�=��{g�{�@�	�dL77q�%�-w<�V}�Ba�Q�P&ce������7��J��e�8�Q����꾨�J�0�2@3I����dH�%�WB�;���{���Q
@;F�I��_���uSh	�Ʋ��֓§�{�2*���kAD�,EZ�J��\��g�o��ϸ��M�3�A�L�xMb�!��l���]��{�PM�xj������#&h����h���x��'���F�I�!r�H�Y+T�>�>�����ڿJUV���R��}΅�aQ�zS^'�Mc�h_��Ǳ�n#R���7Q�|�C��շ
���3߆�,B!�����T��k~���y=pO,X/�=�*~��k��	��\Y�b/M�L4e�)6twP�����Z������H|�;q�a�J�2�w8[����5�ނ��	�����ͯ?���K`-����l��C�{�bq�4�)�J'�0ixdD6j���b�*#G<F�k�z�Su�&s���&�����p5��׉�&_�^�j=��ƺ�d���8�^�U`aUEKR���fh��E�6���8�I����O�a�,T�W�e�p�z@��X�+�A�$�f+��x��������x#�zg�T�`�\,�	�Ԧf��b�g��d�Kj��){}�xK���,��$OZ�1�`-8��lّa��c�N����S������kMju���#ۇ�."7M���,[J�s��:<(F�=gQ.F6�:�|����������x����+�p�K�鯯�˛j����e��K�b��c�#����3�U�2���i�TG�5/!�aL�tt���UG����H"�A�ss�J�D�)�1$����\�
���f�N�v])bI���%t��'RP��8e�y��V�^QB��G
��0q��a���v��̵U��@
�ZCwb�����&�v���9�� F��0 agU��Sp��H��^�8G&��'!�
��2��R��SG���2�c�	d�0��,^;��R��D
wnP~&�.�\j0'�]EZ��l�M����gF�Z�*�AD
$�^�L�׳d[�̚���>��G�D�w��Wx�Oc�%O��g�پ�=þ�F��Fe��*�gG|�7ᐽ�`�<J�|D
�Ƚ����������Qi�壈X��>YF���㮱ϼ�©]�#HOD*�2����|���G�ΒTݾ�'��;y���G^�׽��Y�mµ�k��D��l��U@Ϣb�1�SG�ZB�4�fyҨ�}w�N{+�7�6�!g��M��	�c=��Krյ�+"�g__Q��H�xgb�"�E[��ˑ��Z��
֚I��a������]A`k+���N6I�� y����4�lP�(������s%�\q@���c�=��1�]���@���Hs ��~���p9��΂��~��&c�]����v�� ��%�h��u�8BC@2fM�f���N��G��XN�/�����xZ�(1��;����E�������t7���^T�-,_:�3���׎2ƒ�~���{�\y���6=� 1$�6�B"�2uZ_�����L�F�b�&���[�!��,,��QC%[��f+�)ע8y+0�:���80m� S<˥Kf�:0�FdeԠ����1d1dE��Dij]S��L�<��$�,�Z������д�Ccr=�K&�g����cu4��x'�Q��a�ͥ�4])o�.�����1=��79w�01k�u��9��{�w.��7�'y��v�'?�.�f�e�XCB��wq=n��)�@&[@qdD���yiBc[J��E�R�P��,���-��J��L6y�,:P�'J;�d`g��>w�i8���B�Wk ���$��_���/lCG�_m,[6o8�@|�=�c��*?����?�^}u
�o�Y��p��b�i�^���ÿ��G7��� ��I���yX��H��mK�U|��?��Y�Xd)'`Ң�!���2�����Gr�~;�u4P"�	Ub�%��E��T��42n�ۑ�:ޫc��#8x�ݰlɨ�>6��'��ƍ1o,�_���b �� ���u��/���e;��O�#4�4C�-���7�t^s����g?�%��5���wn��QpB�H1����0<<�f���RMj��,XPD���~�u���Ս[�6|�ݗ�+��3�͗N�U� ��Z�沫09�?�ᷱz�T����W6\|9yzZ�:L�� �L�C��J [,�X��<��tn�>Y7�*�����v����,s�*������+���`܇�'�Ub<:�3t�#��ZOR�����K'�1��f�,c��i��x��OƩ��Qv����U�����ʿ�Pe��ϵ��և6��͢��I�AS)H��H��;�NL�U�jBT(ۙʢ�9e2)�{�č��}�Z�5aL�R�BW�1�B�ז�R�Sro90u)o��C�x�!FH1��,�����Gq��aƴg}���q�*���D������J�bn����[q�Wa�����J'J��\����K��T=�΀}���_'����0m�Z5c %�T
�C�H�D=�L��OI�U?����Y����]��ʈ;8 ��� �Nh ��ҟ+����v��v�%O���A�3�R��g<�Rr�UYֺ��u	h¥�p9:��Z�K�#�
��~Q#"��FY
g<�#7�2[��D�BȨ8I�z�۬��Bz�h~�W�aj���=���Mg,��֯ہSG`��^Ƞ�+T�Hϯ;�=�4`�g �C!�0�16r�D��z�<�y�__H%z���o�v�V>���f�rQ�m��V�=��ͥ�	�(դ��I�=�@�K�=���'��t�!�T>C�;z�wi�W�U�;��]���x#�}�	�!.S� zj
���͸��P�$�O�O�L�$��+��3��<~J�{H�]�ѹ�T�� �400T���%�n>$���������.��!�ˣ5@-�(��q��1H[�o�P�L�VڌAs�)��=o��^��OK� 
{&<x�}�{�]�ko{�D���ق�sĤi]�-�1}�z����    IDAT�?r���5m3�zt��ݲ��kZ/������`ά9�Ѫ�=0=�,VZWd$G_/,2DK_��ؗ(PTŔ���Ҳٯ��7�Y����#�G�_���1@�N*�� �����aK���^}� �2�����i��K_��d��U�}$�u�0���bn>�D��V��:�+E�ԗ��mnl�R����n?&m:�g�z�&xaä|��X�*�]K���K�����(3�(��i��H@�"�_�������>	'B���8��G�0&	Q$�������Q�w	L�t� S��p��*�82�Rm�j6�|H�P$�r��f�i~��T���"�#��]��<=#>\Q��Q�UПg�H�p�+��p�ɇ^_���cj�%�iFJ@/�q�B�L��RI�1U�-���z�8z���'Oê�*��v��(0��w�?]��=w��z�k�@��xnK]r=n�S�\~�s��j� S"	����h.U�����M44P=m�>�%J�V�X�X	��� $@ۿ{���w�)�������x��)qy���s8d�Ux�)Gb�e��W�u�V<��Q�r�ذa�
C�_�m`��98��`�5{`�]w��i����}f���ټ<> u�����lJ��F�:%���]iu�i'�T��r�	e�|MV\������S�7eՔys��Og;���X����\��B�}�ZXu�����N����!)Ơ� n��|��� �M����62�����hb�����+���]v�g?q����r��x��o_|	n��nr�~��g>�y#f��c�x_���x�u8䠃q��a��������m�Z��.�7n�[�|2N:�5()U ^ް�y��1�m{�_���X:/-rR��n��~\���0=1�_�m,�!�|;����.��'6��J������ʠ�@�<�#E	<�Χ�#O!M�n�7d�����N/N��2�g�L�I�%��-L��Y������G�+�9����NOa3�R9-��$�=Z5�a7	t�8d�x�ɇ�ģV���	�����.3�c5|���L���A<���~fʩ��Ǵ��<�=]k�69�N�*A���x1�G�H�k㊨��܇���D�fBd;�z����o����sp�^W��R4���8�����1m0%N�&�����-��oW�G�k�]r`"A�h��\�*�7��ұ8����x��K�̀���N7M���^\v�}�:=@nx��{�y�RiU�P+������A5�@Q� ������A�9����ƘP���2��L���1��v�U����jzHJ���  U�"bA�q�af�(��bqPP���*�#%��@z��}���o�r�yљ�G�Kxy��{�������kS`�ǆ��&�u"����W�u$�Ya�cٔT`��c{�ϸK[]TJ5Ty�ɦ�I�ȁ�H{�9F#��=�Z|.������kޭ��Ri��w{|��B���^�O�D�>Abh?(@�����7Kl,ITF������B�+�lN|��C�����L�h߻&���VO#ł���/LL��@9�d��Po��t����&�\QrM� ?�	�gӐ��=�gi&n��9��GS����')��J<tdU�sK�ӂ|��a�����#�^�(5��x���0�.߄ZGe�-�M!�x�����2�`zؽwŇ��Q���RLT��D�z��M!���u]�-��י'B��'�w���?�k��aO��(�wRm�sn�����N��0Z�	t�%�g�8���p�c��P�"�<� �~��X�6����Ǎw=�Zl ��ԩ��Rա*�;�F/������*����Ӥ��N}Uغ��l[F�L ��[�y�\{�����Q0I�V'�=u����۰��Y7]?�/t�^��B'fǦN�i����A�Eg����8�cx�a��2���V���p�qּ��b#�<���ͥSC�]E�RBc|�j�ʨ8C�5ϜT
i�3�ͱxA�>���5$�w�Z;�d��3-�Y�@�I]'e�̟��H��b`�<Ē4_M!�#�jEo��}��Q�J��V��m��#���80C;9�#���b�:cJ���(H���2�)o���8ۖ*hs� ��T�ٺ�E7̈́N[���`�M�5��Q�`rl\BEm���<b�8��q����<��I����S�;��C�3Ti��*'�]�15+)�+a��?��:d۔��ķ��8����ݥ�榚���r��r��\��:�D��V�A)����}*�vD�U蕪�ȴ�qtꤟ��e�P�F���
��*�'�8��;
LU�bM��:b�*R�
2ſ~���S�)��ο��9�T&'ҳl&���y,�7��b�c��n�Z,s��JYK:�&ڱ&����s1s�|`��I�m��I!S(H�B��*��� ���U�x`�5LVSb��b%�zI2"�՚�Y!�ZV�Vm� ����E�m#mI�h�4�zu�F�:���8�Q\���C���p^E�ÓO/ŏ/��05��x�	54�w������o�v�n�o������1�c�h��Wx���vǏ�u�����X����
��e�i��=���F�) \��K���W�\�Ѓv��k��~��7�{�Ì�^|�����[��8n��!�z�=�Ǖ���<$Ս���7����~�7ޮ`���4�W�mqN�Е�P@����MW�J�&F\4�
�y��
KMQB�<r�H��=@dqʋ&0��Z��FI��Ao���$ɿ+,A��vi�"�6G^��g�QC���[���2��É���v�[���zia�*��*�b@#�0^{i�t�SX=�A3Ճn:�&��H�8#��4� '�����1��(�<�3L3h��W�Lɣ"��ͬ�nW���E��: �sA���9�v*&�D�4��1.�#�}�l#��5Q;v�1��a���-}&��J¦�,�^Wɏ2��һV+��S��b���Sp����qPt��=7����U\y�}�8�F*3�f�+@0��i{��
��l�l1��:�����i�\��*V���Vf2�[�J�`��%�)�x��+��dXOd����e��q.l��Lo��{��(LH�/]�y��S�;v�O601�V;d���K����	�$��J��ȳ�r�;C:��ôJ�K�>�=#!`���p��C�T�9�0�e4���%�t�s�ȗ��	�*�����%�+�1�#WeLI&�"���+!\f��6\b����3Es�0y6�3b����.הJ�*��T9����{z�s��A��XrK�����+x��}iL�������<��7W@)�>�����㉨���}t�x�X;�|��"9t���/*�~K�7�ﺥ\Z�
�U�"�'���� C����N/&�¤�x;�SEfuʌ�8%9�"�V�ߴX�E't&����g��]��d	��$2�*��ׇϞ|�����E�b���+8���o|7��,�O���449�}�i�}%�!��+,J�g��)�Ӟ	JE�S�*A/��U5�]%6�\x)�H'��'�y^D1fZc�}O��I��_+�La'mOGr5N�iQF4���Qa�T�H���~>����������?�V~]��å���K�`"�$a��^����	�zE�w�NpZF�4�Zi��*@��1I�i�� ����I$2L���{���sT�͎�+D��X�"k2A�L�Ҕ,�C��V�gz����X6)�RI�)�V�>3��b�h@�90ur)���ZcD�A4O�}.���$���<:ɤ���J_���1%c�����Gc�h���bq+M�2��0��I�4QI�N�@�d\�i}���S?��c�Bm��$�f��1��"KƔ�7�6ʛՕ��C
��,��[�1��Iy٧ʼC�Bd��Jy�4?j�%&����i�[G��[���${,�F����V��(�}}CC���Ш*cZ��4�b��e��Ho��eD�P�6�V��̓��@��	��xqq�1ù_������ى�s�|i�:�,[>$��,|1�`.��|�_��6ȜJ��YV@�T&ю���,��f�w6j�<��d�jN���TDv���*kVA� Vt-Ib������8�+�ψ����\p\��Z]�	�����˫M�D�T
�VC4�AH�s�6!6��Ŝ��55d�p�c���?�����v;Mڤ�'����"�K~�=v],ۇ�F'��n�7�~��;���?#O�#?����
������_�®;�|�l��V�ilu�}O��+�F��Ƨ?y
�<����V!���*��c�˯�K_�>��} IA���݋���������G?r�H�x�T]\{�=�����$��/��ٽYى���S���K�k64ЊeHs�n�����e��L�19YC�Ά�HS	��Ez�����]Z)�D�#��:��m�l���33$a0<��	`�_ �Eg_���%񐤒UoM&R�e曵��0(�	���A�E���,̛�=�X�]�,�V3ѓ�3���Ē@�����K�����Ͻ��W�(̜�D���suY����2��[��:2����v��zf"VȠ�>�.�%�szc������� �F��h�1mŒ(LDq�4�S�@��j��j����H�֚h�Ӛ^�$�Bc4�gØ<�G�%��p�����]ֹ|�.��q�mD�1������7>��g>(R&C� �g þ�t����5`�hVL����Y��TZ��UW�'ɶf�R��IL�Z*}��|X���-;$�E�
�|&�; &p��1dB`� |1���D�㝲<�h�)��w�I4۔�2&hU?�e�!�V��I)jR@7d�7{~�~˜ؐi䬖l:W��ʀ�8��o�n��3B�lɘz���l��Rס�+}ށ���Uy��,V�r ,�k�����i@B��T��hB�}�^���燆��Ə���6�l˽sp�j�W��4��7����Jp9
��6�S��zv�H���� �g��n$}�.A�^wMW�%N8"��kN*z�3e��Q��㋧��:n���#i1�	c,�JxeUW�� z�L��ht2H��G*�F�܊(�l��Tˌ�z���<A�<�8bp�
\�p���Z��ǹE����2fz/�����f�D��d 0`]-6�+��Tq�׹�
�C��_�D�^�@�6�����	|��Ǐ� �NK����UIe��~d-~~�=X?�D=�C'��d]�$�#N�\[�^��(c*�Mv�8�d#kŋAE?|TƁ�<�"˹l�B-��2.+��/c8i!�����g���6ޔx�&�[;4�E����KUA���]�-�J+�;�����g_X�P$>H~k�'QI�R$�����F]TEu�+2�,�-�{-�QD�gЫ&���c��X��f���H��G��������X�R��h�ب�7��.��`�gc�^T'�x���x����8�E+=�
*���1A:��|ZNq�6s+�?kGG��Z֟�:	��/G2��n�����'��)/�*��<��i����'u�T#Ҍ1.�bȘ&�9��s�5�I�GPK�4����^52ڰ]����[�F��LA���
L�CchL��m2�N N5'�l��Ҥ�z�jA�w��V�g)��f�}{ݖb����r\����W��	���n��1	d��@����u L�ol����% ��br�=��樐6��o�򘽨���ԡ�ˀ�l �׳�X�~�[D*aݎ��8ȚN0=�'�#��)����Χ���[���0��z]d�s����w�E��Do/���h4�,M����|��j�.�_���J�e���CO���;�G��k��WYg2��Wp�z��u���/�����&fރtž^d�9�~9�-�d�.g��O�ڱ�!#5��MzMd(�iU0oFo=�`Ό~�`��>�^~�Y������H�8f��p�O.����o|GuHPK+㺛nÃ�<�l.����E,�n���tcX�r~t�O��3Â�[�{����}�<�~w����{�!�ԓq���Ɠ϶�V�5�����x�-|��c�SO@>k3��1��7W��;���.;����Sy��r�]~�H�ٯp����=w[,R_J����a�隻02�E,݋J��\O�����K�g2��3Pٙ9R�cx��X�hR˴�!G��2WzDA�$~v���U)lM�Z��b}o���_�L5��	�g{*j�����%�,$UQ�7�t9�g��Q�''��Ԑ���, ������1�����~NA���c�xs��l��D�N5�?韁x��L��i-)�v�P��Q�ZC�R��((d�1��b?DӲOl��Vjh���?5�l���2(̘���Aq����x�d�*�`ZF��n-��l���	0`k�w�%��7��v�H'�2�od�Z�˛�pN?����;g#'��jtP*7��(�iE�6��=�2���Q,_9�n,�޾�t)4N�9����X���gNm��[��D�K�"���9��I����Z�w���{��*�N�Y�qV���n.�D!�n:�%��`%h��Z��	LS��$�� �z��=�֢hPHZ�������5�H x�t �������0��p��-d���' �!cc��1���r {u]��
 �ב֮l	�q/����X�+J�|90�1�g�=��b����,�V����Y�&��^�_�1�S��Z1.+���ߙ���qYG�kj#c<�ykD��)y����~]0�:=i��l}���^�m����|�9y�^ �E����+�����/���z�t�d���B����
H�z>j0�2� r[��
�N�<��:-�3_��m9o��M�����:0��#x�z6U���=���)�օ���B���P��4KC�6q�A{�S'���b�"�J�S(�m �޻�^�U��f��90~��-3c�bS��E�^���F�;���� �� ����G�E���L4oFG^���������%M?�޾��
U��"���<0���[�C���O8BvQ��6D�زV��\ό0H�kN�.A�"�� ��@�s7z�� U2�-��l�Y�<�2��q�ce�����S���y���-3Z��(�{���_�j��U�;�t�0g�~�5��UF���p�)�c��S�?i���]:��zO,]��FZ\�鮔�DY�d��/Oh=�b�bIuڶo��{$hSYe1?�t%!c���"�i"0����CfiJ���F��q�FJ�c��J����d-M�Ư�������R�
�$�L��$�ʙ���K����k� OBQT`]��$��y�ͣ�r�4Z��˳�=��,[l]	Y�%4K�H�!���_��T�mW�n�}Kf༳>�g����z��m".���*�|�cr�v�q+|�����^ۈ�����5\��{q�/�Q��3��i�r��r���=d�VaK5�����2�O�ݴ3NV9�H�%n�����8�9�x�x�;C`
੗F���`J�3�z��h�9��C^�.Hk�0��lqy.��+�vx��*.���X=�A$��Y�(�e?4GG\]�$̩W�E�k�֥r�.��"�6k3y�T�xY�fo�c�9�"��!�~v�5&�Ϯ���1P��'Ϥ���������p�!��#G�G�,|^�.��%���{���?�����:��f�f���?a�+�J�y�)���r[ΐ}�)��W���5���ۃ=����������~y{�i��O8��!$�:/���O.�����6c�=v����W���������^{}���}��y�bۭ��6<Z�w�^{�MT�e|������,�[��q��7�qFǚ����R� E�z��X��6�i��P,�؅�u�5�~�SX�j���)
�Y�r!��{f�J��9Sj�-�J]`l�'�'zB���X���{�!B$A&G�➠�!����;�L�X��1�m@�^����w��    IDAT�SĶ�ؓdJ=��G�y�F��X�a%�K�;����a�N�1o��H��b�����G�@�5k�g���=����-�QG�T�Cрi��FT�lI�%�/��j�\���:�������H�g��gO�Li����"�d[�b��0��Zq�85���[@��9�da�4	��&8t_��4��эk�,m�[��o	�ݵ_��|���<�䋘>}:޵�6"a瞣$��H�?����^^�	�X�1ʔ2�r�n�`tErD�j�!U��P7o��f)���23&�2~'���`�b]I�Y��+�Q4��3N�4`P7!&e��QU<�C��"����d�VG%L��NC�2�j�
ʬn�Y�z�������\���5t��#����l���_er�" �.�U��ZD�E��l?�mv���J�d�s@#�ZGf����q��\������RAs$�3��`�G�%���ߧ:r�)��$`=�:� *D:��+�Dr5e�5�5�lD�,�_eZ��#Mn���n�����}S�����4�q���A8�&�XW�3"��pvi\�mX�]����瞆���!)D��2���lϿZ��܋'_\���O�jA��4:r&^<-���1"S�D��J&9�1%�����O�^�~=���U���E6{����5�p�S�4�ת*.X�9e�	���k�N�"�bRĲ�¥�҃*�����u�u�J�hW�ї��}��ӏǎ[%��s-��P�=_���xi�$��>tx�Df����b3��Ŷo�5�lt�H�K�+ɖ��!3Ί�F�w��z�4,�����-��=�D�tP:���b��4��Y���~(��p �&�62�S��>�}�@�@1���#�LI�%0uP�om��`|��F�R�B���L�.�iT�q�|���
��	̛��>�nl77-E�����\x��	���b�X�x��W���"�<�5�h�6��#ށ�?{��<J�U"	|�YZ¯��O�����Qj�)#��	c����'k��/ވ(UB�=�*��0�"�MIi�\yE�
����x\�)qkc��6Li��@�JM�y�ӈѡW��;J�80��7��cy�$�b#9��I]�4�4w`i}�5�N&�7)oeӰ0�$���;TfF
X^(�vȘ S*�H>����*S��K56k�)��N�s�͏�]cLǀ����㾧��h.�r�I8��5PG�7Vŕ����G�GO�td{{K�L��)6"C��������|��'`�qy7�����3�<9�@ݠyO��X{B��ٟ;?n?1��r�ᳯL����U�b����+����3��8�X�V f�)��hg�W��Qn��m|�����0Pi�gs0u��t R�AȬP�.��j�W�Tr�r,�W��g"�=�*���s�lVd�d���,��{��S0��b���fi4�lOb��f᝻n��)t�U�
���Ǟ��//��s���c����¶�]���ַ�v�f���˒������^ؗ^\���|6l�$�j��;����6`|l7�t+n��f����:�m��\�
����v�F	����<�3k�$حVW]u#���z	6���o��w\,���+�?�	J��pp*�c���:�0Id�����������g~6m �Ɋ�"���S(M�Q�4����X�\N���c	�<���n�^)Z�"4Z�z�-���0D��M�"g��8����B��bm��
+����Țe�23�+�t��� ��7�W@�A�rpmpoH_�1|z`h���F�|�M�-y/��$�'F�q͛�wq�ߍc�sgdDY &;-`|��MC�X�����7�'�Gs�.}�~|ዟ��m{��k���.ǽϬ�d7����쫠#/�^�-���i�.[H�,zfJ3>D��0C0�Lu\m���+�g��e��$�3�#7s�L��e�=��}|k��'�c�-1P����y��a�Kc�1�~U���(����J����[(QٸNzLo݃�;��܃LL��[���JL��8�S'�}wF�ى�-`��{d)}j�|{�nZf3&��D�+�ߦ�4w^=P�/ɲMg�D�kRz=,� �M��	�n8�B�f�N&Ҥ�$6ٳ3>1!��dL�@1J�H��dZ~���=R�E��xK��Ѷ�(䋲��8�[�z�� ����z΅U��{L�xmʘ��WMf�n��{�o�D/R�q���j�5S���8#$:�$F�EuՏ��T�</�[�)R,+�^� c[��8
�lA�a�}��J�C�*�\O��dѨ���+�#�]L��{b��P�O�4��e�A+��R�kKj�TbY}��P�]��	e���	3ɚ��߁�+E8�.ޮad�r�4��z�q�ϙ(�Ta�=Ǣ�=���;|o�.���E��@"�Y)�0��^�I&�U�8`<DBn�[~�7$����l�J U	��̇�����k�3�zFi�'*.ϱ%�g-š�1���!��֧l{�_Fpf�f?#�NK��߉����Zjp�n�:1�nc�x{,���}��m�L��g�X��g=��5����Ͻ1�*�⎯��ڞ#���x�y(�uP��C�@!�J6���۩(�k����޺(:�S8X�fDh�=V�3S.{?�s�y�9�f��!����0�DUW�قk��q��@��5E������$&���΢G�N�bN����b,#��l/Kw+ȣ�S�?'�.�聸9�9o��6��p�3��w`�h�d12�4��dg��&��h7���큯�y�g�v���t���"������oǲ�c��XT�!�a�ɤ�R4��1�Q�9�:�ʭ���ow����6W�4Y�e~OykOq��ӿ��C%�ku�4ۢ��(��eZ檏!�R*��S���3V��bFP�-�!c��2�CӌӔS5a⽔9�dk#���y��~��P��v�aVl���s���ʔ ��u�YF�=��v�y_9;�ɘy��J�.�X��i�1�5���?��������vs�ϝ��޽�&jH��M\��;q�}ϡYO�pR==B��h�V�J�JE={Y砉���I�	��Fcz�c�C*�9-�������С�,����g?�O�����ʺ���Fq�^�WW���D�VCO�,������w��2�c(X����_�^X�8�+<�z���+�jCS�i�Liqξ�����?�A�L8�<.A����잸d1�L����h���	��9�B@>%�&A ���K<�QG1��¹��v��ȥb(�s�ʷW�4>�����4�z������5k�ꭷ��J:~��Y���C� V��#��buDp������v����駟���z�z��S�J�F�81��Zk ��ϛ���,�822�xc�RB!s������Ao?��!�z{��$������0g�L�{�x�ŗ0�a��z
=�k;�,��������h%�/@ήb_ao.���={�Ω������o��3/�C���8���O�D>-�@��@V�i'��/�B�b�tZ@9�8?�d�/�N �9Q�8��G��*]���z쬗�*3V+�n����fL���}�����<	{�ԣc�� X�%��]�ѧ��/~}%�|�%9.���3pک�bz�9j �=��>�:F�9�)�O��e�.�唚��&�(o`*Ά�<zgMS)o��M��r�DHj���W�h�m�d�l�Vk�qUq��f�0�9����[�(rw�U�M�qJy�t	�d���%�  N��S������޺�J9'�V����f4+C"a�����}������yx).�͵ذa�l� _<�cx�s�CU��y���Ɓ���>��/��Ϊ�������u�J�����5$)�=3�e�?-��I�{.Y��%	�*�k��_ m<�&�<\�6��FQ�W���Z�a����a���\u~�1�]�`�]��d�c���.av=)s�d�:�:���;9'�d��I*uf���)�i����F�BPr��%k�� ��2�ia ��B����`,��fV"�iv��{\��C<��h#��5��+v7r��ɊQv>[��LL&�~.lc�{�.�Z �D9�QA�c�(0����IF����ȯ�g�>F�g5�g%�$�&G֢��=�n��fO�G�V�[����+���5�4���"p����#gp�xb�e��h�a�ԇ��GE:Z��_����]k`��%z�����)nr�c�Fz���E5�Z����;Pf���O�9J���bM��F˪���j��M �Z�q$�%���e�,|����=�����8B��g'��n�����_�̴�LQ:ڊ66�8Z@��-(�;��Y�V��~��l�RS�f������~��^ :#�4	��'�'pl��=s�)|M˚��a�
�_v�����b���y��=����4�1�����E��`�[�4W�*�)�Ϸ���t�K��U�b�8�]���_8[O� ��(�����ʛ��]���-$�E-�:-�4؎W-�Y�>������	�8�S�N�g�X8R𱿍�'��o�� �^q��ХW*_2�A
#�z`�F5+(�:
n�I��7'��L�g���E�FCM�c`&�+
HY�t�;*�M�"�S�[�̷�ڸ�-����Lʛ��ソ��)�!�ψ�W��d�l����FI$��1F���h~D��3P��E;R$��S
�:b�J
��iAS�utZedZ#�w�|��tn���ֺݮ�yο�O��g�f,�f���p�{0�#�����ww��{�A��@��l�Y��B�i6Ԟ�I]�5�;-��u�oV`�C�	~6/�< h��q3�lV*"Zu��& X�vj�w�HvF����O��`~�kxj����x��	�A���n3���.�drI:r֑�aoZ�>m@�f���.�rs����� s]��Y����H�d}.;�yw�6�%�~�	Q�UJ�c��&�ڻ��e�u��˾S�3%G�C��	j�9̖��Hwj�&Zr@3,�S
��!�-�.�Z��'�:�Ceud7���	�k���V]�d3���'+Dd�)�i�o2��na:;�Xk�[C6 d�y�\ɄH�EZm3��,�|M��:�S�A��E�C�M"(�6hnTo#�̉ϒK��\pS����:���8H~��fHE9�8�F����.��gA�t�?=W¹c�bZ� =H�f�0����B!���������`xx�h�!�f��{P�Ʉ�,�U��SM� ��cEx�;-qS,�oFO��ϟ| N<boL/�D��%)	J�U�����%��3�\���5��%ZO �m���_�Uy#�^L����4��O��$��56�C�K�1��\����]yY\`Mb�j��5��n�Re5����L�C+�נ�T|�]��Ĭ��i�%�hMLJ�i���Ȓ`\L�jPs���J��;X/D�ۨ�\C�2��3���g��A�Z��"0V��H���04TF>���.u���s�V�&s	�l ?9�?_w?�xc&�'�jMb�/�i=�f�b�DP�C�%lʼO׼.d�q.0U�N�:���H�2�I�qM�68\N���\��24��#	���d?t�-.�f �z�Ȣ2B^��UE�XVei)���f�[˪_����j¦̟��4�hҢ�Te�
�k����ˣ�l��ag7����pf�3�S�S?&��C.�%`HM��
Otm�XRml�\K��$�~��O)G�=.���)Z�����������`�����ɶ���=�����SBNpw.%�mn���R8��a:�?���r�@��}��!0U�}oj��_Dk��R�I�q�y�u��r�${�{d6)�U���-)tHG��UU�s����Qn9�t��<ڊ1A�B��8Q`�VA����r��ۤ��[ly�)$<������)�4 ^�"I���7�`����Z��2�j�(r{�����D��{�D�Cbb��$2�*�M����#9 �b$V�v�����gV`�A/�/�9�x���X��W��Om�jF'kK�J^/��J�ۄE�J�l��w���}�Kd��GGaq�L�g�{f���[����o�ʠ��#1�Ն��
g�C��[��G���ev�#�
}D�.ѾY���K%W7�3�w�1��Em��m|��p��[K��]�^.�S6��[�	W��46�b�&�DUB~p�$q�M�*��Ma��4�8�p��ŘQԜF[r,|Lԁ+oz���nT���؛eϦ�U)y���'c�t�l����[w-7��3�z^P@@�FScL�4t���b�B[���Ḙ�L�ę�f�b;�Nɨْב->�E= T=��Ǒ�|qN٘d�7.�4|��L������^ˬa1����I&��H�F���2����4�pj� ~ 
Lö&im`�ǼXp:��l�q�i��ͮ���o�A|�˧b����]�K`������_\�;xF�n�`_:�q��H�Uʻrs����g�i&��;�x��P����nRe$�u�,b�>̦{f��j��ѱV���mT�1$R=���4S@�Zs����D7^��j��D�E[�I�g�v8>y�Ru�/V �\6�o��:���3�a`c�SƴB=i��UdW!C���F�����g~�4̚ѯs��������/�9�Xv���p��.&�J�($�ْ�fX�{۰������V	�-I�i�ZLH�ْH�=�tȣ_Y�C�޲�����,V��5d�m&�s���U� �k�++�L��&j��dB��| ��sM����M�S�L6k�ZgK�iڌ+&�\�4b1&��s���G7ܴ��c$>i��bF��Et-����5[˽�����8b��b�a!cO@��8έecw�t��7�9�l5M��L7����W�p�3h�i�ľߤ0��_*j�DY@��!�\	q���J%P�-����F0�Q���2::��RY9�5���~=�������j�#V�m���2@oz;.(��sO������R1)y�j���ѕ:��+����e��ރ�s{DzBvu�\w��������,`�ҏT�,�m�wH�m���hI͏x�=yf��J����tP�٩Յ�lU�c(��$�(N���_�������NU��N�ǴF)�0���0��?�P���Redz�G�nj�cG�/�k��ry��0P���C�������N
��e����z�0���ɧ�h�\|��c�������t�4��gq��ϠUn!�mb��f��vǢm�"�M��$��TԪ�r�v��񀫷0Yib�h��؈'�{o�wB:a�m �F^;|%��cU�F��l��i=Iq�;���m�/��WU9~�wu�%�f�����Rkb�\�����oㅗW�/J�7o�$&�[�+n����9}fL%�X�Ģ�W]�C��	�zb���vS�I��W׽�HBK �:�F��&�.M��ޘ �:SeD�$���&�¢�DT.��#�L�tN�"gr�P��]#Z�O�+hO�2��
��ْ3��!���FV@�$*~�X�4��./G�P��>�/��^�:\����\I��Y�!#ղ�Z=����%�J�L�Ǟ�L�KuU�b����-
(�Q9o�`� ����:�i�B$�����d+Bz/��Y�����������Q}������=�R�P�����=N��*��jo����x�1�g,���hpnl��N�#�*�%��m��v��t/��
O/{�x�i
r���Y��a��EרW\��)�Ȗ���)R^�q���S�C����qe�m�6(��"'(�l���0`1؟�/(to�uo���W�����QE�>��(�Y�+�'K�?�����M�<�܀}�2�lq���<.����LeK�S�/fg\�tl���q��Oas)��z�lN�'�b ٓJp��n�Z�	#K���[���ߋ#޿���r�ŋX�n�&�/}��x��:�D��雤���I�b��9bn���g���)�Bl^��5�2-���Hy*�e䱞    IDAT��`$����b�w�2.��yDrI���u�-d`*flR�:�#�J I6�\A�SG��(&�4N��BZ昒�᧦z��^��t�%n�@)/s.�R�+�ԅ���R\�QDJ�vL��3f,�w[���+��?���ʁ��)#Z^ԥkt�ݚ�_^��xN�����O���Ƙ��⧗݆;�}�z�}��<��$-��:),�f6=��x�޻b�t�7��A�|�
��j�>�<z�9�X=�j��o�df�j��	��wd	j�	$�5$:����ę�>,��b�KGp�E�a��
�M�i�)-�*c߸�V�GNԐ�u�����v^���ι�n��Re��6�CϮ�.�olh�ϣ����Rs���$��o��-�o���YUf1�nMܼ>;)4Y�o�vS�Ȍ?3�6Zؑ���j��rC�gC�8�VYg���
Z�X}��c���|̄�������:��#$N܈C�|&�c�(e�������_R^����ֿG�-�Y��gE�)�<3��5��T -@ҿzZT�JP̿���J�K�R��5�T ��N�	d5��{��F����ެ!o�쯜�c�:(��o� ~���p˽/���#���G D*�j��S,eK��	~�"��3T8sˑ:Xگ�V��F &��&���IY#�^�|J�_���v��MO6y@�P]��v��������`r��P�����k�v�Z�gϟ;[\�����8��/G���V݆����w���v�4�H��N'��-�j	0�LT��y����䑟ޏX/]yM��� �{M�cZ��J��p�3�#?�-S�Ѡ,���-���Ƙr�͏Le���� ��Y���RA;��le=�հ'�z��ju��r��f���>�hk̞7Cc5���06m��oO����!�zR8`��qྋ1�?#���_�sˆ�q�$Z�%��w��ӎ�.;d�����t��_�P�L׀2��j�X��c���C��C,���QQ�2P6����f��#�j�����3��~�Dr1����4���u�m����/��<������x�	rX���x�#�`ʍ�t�� �di,VQ���ǣ	Z��¹�!�f`2�fI8�b�3�IB2���>>$L�6рs4�T �E���h�AEz�� E��'�f8��G:���91"��{e���H����s�V�a�/U������>��{Yc���]�ȝ�:`��^#0Z
At���s;>l/c�'ز���:������PB��Yd�~F��М�+3�R5�z���1uQ#U8�m��y��J�,��e�+���,�sK��i�;އ8��˽���K��%B>��������R�`-Di>�!S�\r>S:��hqC�=Yd9�[��86��F����aYUV2��ٔ�\b��)�s�y��Hn#�74r����䌼�?oA�i�"��n� ��qW�����;��_r�"g����I��ck_kh�+E^4d4m�G���1�y�񴿌��G��Zd�'��kL�V�^g��y�v~�J(�1�~~m}Ss�0~D>׵���{��U��:�
:�1�����?��E�h_$�O��]\~�����o��D�*�Hu�?+�bq'�+��z��Q�G�`n�>�s������5ZHb�M���q����NMC"� Iƞg���ΘjX�Mj��C�����MCLB`*��=dL�J]��$��$�@��b�-T�G�/�]'0�!��t�$8�o�8cMP ��!G ���Ą��(女n>�T�+ 2����a��iD��1 ���*�����fX��р���cA}s�>��]yS�!�� ���'�d^�gL	L��~{��__�;�{�F�g������	4ANn��*~r�͸��g�x���/�Vc�`�=�ȃ߃w�#z�y���[ ��m;B��oWp�]��G_��5�Hf������qA��Je��ӏw �v�q�����_���.�+6T�?m��(bPlL����-�6&o�'�/���yx�p��sgH�O$�H��F�݈͟�ֲ�ҋ&�}^z�Y�R��|�^��;J�t8�~���':v ���W�Țri�|A�1&�t@V�۪k��T��3q&�L��,�82i׀�ܢ�/J9�_���`
�l��Sb+��jdFd�PR��H +�U{��:�t��҄M��xx/êYC7�R�������Y��_� ��I�(���;d�����*͔��I8z�٪s~��׿�%�;`���a��ރG�Y�z;���݌��k�Z�1#�~]$��z�*J�i��L+�A[��T @���w�פs�0����@��RA��%���l�-��k�U��F�1�ziN8�]����A�R�8PoO=�:~���b�k�c��m���~��+����F��Te���w����<���H�u�Y�v�v��
�%�'J�̓�����[L��^�`ԁZ�h5�n��%4(-i�Qg%1�Fa�4f����g�txv�ҝs���)��n	L�Ƥ���e���)�c?���1&&p|�J�Rݏi�P��P�EmrITQHױ����������Yl^zi5��a���
�S���p�!�a����{j�6�C_8���O���^U���lyX	,�,#���k-������z��1\��Ѵ����J�,�N��@�QAO���~��8��c�M��:����ʣ:�oa�L�dj���7q�ewc�Ɩ����dKu.��� �r��SW�� �X���[�'�*�}<���`�B�T	�6��c:ר.�_��:e�K�@}aIl�0��odE��}Jg��D�a$L����/)ۡ��z�Tj�pP1gX��ٓ��G���%�=��T���&[�~-S�tO�#��_3 `ƊF4%z���Ղ�~imؒ�� ��^|C  ��qN^�����T��r�c5�BH�*ZT�dϒ|����4�(��=�>���e���,�Fc5�sK�(j3���H<�&<�٢ó�����MD����R�Ϫ�R�I2X����mΡ�U�?�yT<�'�L����d�)9BP�կ����Nu�i��󤪟��+�ؙ�eA�*�����M�t!p߉���&�3����I�p�ǯ�u��yz��?�qg3C��k�Iw��l������w>�3�R<v�PD�o�M���(0�z]&���P��4k�ٻ�d�1 ��"3wY�(#�#��б�Z��B'UxT=u�t�8d�E��9Gcf��R�Dq�j���8.���o�(�D'^@2�sGy.k�?M"u	�A�S&�TQ)��4���8sm|��#�S�D?�6��rI��?=��\���i�g8�!�n"LȐs'�-�8�E�h��`<�|�#L[$%h~�[D��a���6+�F�;q�i��FmxLf���Mm+��*K����&ͥR������V0I`J��?������I��`N/���ؼ	4ɤ���sL-yd}��JY���a�ݧ��{.�f�
4�hREK��1$��w�zv������ǔ��<�Z��y�z�ӏ�q���D�R\���/����$�6
t�Mv0{Z'~��8��}�͜�WPj��e6�9��ъ6��]��K�p͍���g^3�t�_�7f*�����#cb�w���s?!���Ch�ȳ��ݟ_/�iO߀H�ҩ���a�&�Hv�h�'E��jՑˤq���I��m4��[�Lb�	���'q�}/�ڦ�k&0"��˒��$Ҭb��b��&4�� _��[��{[�5	��(A{H��f��j�D6��V��&]�X�R�&bd�YN���N��J����V9�I����ƴg.~>?�OV���i�J�BIP�d� Ήk�u�̫��T ��*���W���8�;�v_����`�*���À� T��<���ՠ�=�54�u�.Z�-���¼�gK�3/O���y5֏��9B �t68�	�7�F� �ji#~$��K�����i��l�Z��LG�k�+�qL'iR��3�9�UZ��B�.5���G�:<j����q'E>�6��	T'������O���s��K\s˃���.��U��S(���g�s�m�l�1a´��F,�a �?�W��*6Tsh0D%ēRA#0eO'���K>�Lo����I��h�;<�$�|����϶ڨ1X��h�4�f��W�R�2��Ԙ:�Z�=ADM���E�,2a����H�m�6����ʨz�k�]��<��*&F7�4�^��;>q�A�q�pt"F�G]�+.�	����b
g}�|�Ľ0m@�+W���#�<�X���|�<��q�ɞU�>)i	�O�%"�&���m��M�Ҍ���[��E�`��MRd��I*!}�<PI�&��F��vm����Y�9G|`;���T��0�s��c4!�B�B!���!�����w���)�r}H�rJ���V��(��і]�88�sV�*���;S�=u���l��ݺ,ij������#�C�^[b��kK\�df"��)9e����M����y��;�S`�̰�-XLy:,q��2҇�F�oDQ�?W��-�ʀ(����vf��:8@i��jb�`�$�p�L���A|�0����`�H��b�Rg����c˘��{9�n.Ѫ���|���*a@Ss+pX?���R��D���<�6��|f���R �j�cgt�d��(MJ��%ڿ���WO��<���lA���,���ҙ,blS��s���elY8$�5%�]!˥�� �E�Ơ���)��&N����1J��>c}"RF��������͹ًS�=� ���Va��n* ��Ra+��A]z.�q�_^?�F� �������?����
?*X�h鹗�;/�h^�Ss8˔��W򄈣�0��>DL���?��5#�
�(i�0�2��[Ȃ�~��z�&�F��Z�!y�������{{]��U�k��W�֢Ɩ�܀�yP�+���P�5*�i#u�f���S�<��kkU�h�☃��w��l=#-�a~l�9�ҫ���<�Z|�l-�Tm�D�'�cv|�XH�e����u[�C�<aʃ�1���7�c�ܣ�d���P�<*s�;�,4Q^[���+������TSW��-S�c�uJb$��)ݏ������=��1�r���:���=�y�)ݷv!-���OS��(0Uo�V��v}���پ�9�SX2��dL;�١K����>�J����{�O���.d�p���M5\���q��"�$������������=��$)�DV]EC!\xB'HJ�(�Z����\~#���y��� ��I��js��8>|�;��o~
y�	H ��s��ݟ^�Uj������c�=�C�.Ƃi��c���)�3m!����?�$���.��Vl.��`�+�Z�Һ��Dd_���E���������h FM����JR<�b�����_h�D�6�'疖Ǉ�i14�M���X�.@��4��˨i�0�[��h��J|`���(�2�ڇ�]����
X9鹁C7J��ʰbeD���bO ����i�4O5�p4G��Z}�5�P��X�[�X�^F�^��S�_����E,Z��k��7=��o|�X:mʐh��QA)���.�Y9iP�Y�2v�&V�Q��4�9_�R��Z���n� SI�h �D76�$�
L]�&����ԁ�&Nd�ix��L��ƉG�sN�=q��ފ���_ǅ?�K_Z�X"�l'w8�8�xl�UNfo�O���]4�1�������]/c�Y�}L�9�'�ɀ�_���9Ǵ���e�{��ևn1%��r�,�{r�=��AJPYB]�vQ�1O:���A�M�/�-}�%J"��uĕ7Vk�<�=�i��������⏬�`��6�)�T٫Mu {��݄��՘�|�s����ED��u�8p�m��K������'�t(�:�(̟��0,���[��{�q�*�x��(N��-�)�@T�pQ�s���S��(8�5�b[��ke���˰n��X��L8ύ�=�E2e���S�`���< �����/��P���Z!2"�YS�P��L�\�Â}v�9�`�w:҅tY�HR���Lp�&�k#cE<6�OI��9�����B�{�g���+aL�|K{v5g
{,5��Oʕ�܊��7��.���O~&H&��8��-v�!;��ipP��(}��[�W6d�H/��x���US��jd�BS���9\�*�^�0��|�~(��rx�䌋�:�"����=�m�<����GԀ�����Ds��ۍ����s,n~��e�9e}�lA�Iq[z��$��Y��ԕ�v����TQ���[H��fM����I^>'c�h*�j6Q�TP��16Q����n�D��Z+��� �b�y�SYp�p���h�G���(${q��N���� �;?�<�������ew/*���M UedRy�\��Jrk���7Q �%(,�>�Sb��� /�BB��}�K>�0�u"��Q�L��i9@Pd�]h�4ڻ~2�$тQD�ENL8��q��a���SS(�����5Z�G������A���:����GsZ�(�W�tiV6����}�0�l*��I,�����?�	o�m��ʢϊw�l��V<�܍��і6�7$j��ѡM(�nF�>������3�pvb��N`Z���^\u���J�D<�#3tc�Z�������J��8>�'R��o��-k���c�����!Ṿ�1�2��uE���dK�qd��W����?�sLe�$Ae�LrVL������`��4M���ҐqB��cdn9&v2nF\�m��/K�<eõj�s-U�ҥ<�[���+/Y_�-�W	�ӱp�v)�|"~$�:�� �w/�÷�zZ L�F�wy���1}c��K�����J�g���O�������-_;��/�����h���чSO8'{0�L��<�h�H��oAX.�/6�z���a�����8RG��}�	-���t�Ht'p�A{�����$|e�}���8�'�`ŚI$�Y�9N������8ffln�������2����/wq��7c�PK�)]rC�m�Es�/�&�2ٝ��y�j�ىȂ�]����Q��J%�0�_�}����Ny��Ko�jI��*��8���5�*���[`a���5���M�R��<�F�'-%�2�S��*����V7���FMD�y�G���
A���-�z��X��2VG��*� ���R��B�@?�����z�NX?R�5�<���H��!�AFN�A*�E���ݏd0�T�*�
]�Y�'@)/$S2��q��z��J�,�T��q�2Y�sYE�l�Q�Ͷ���>f]#�o��ƚ�^�vJ�9�ݞ���Z,Y؋��SX0G&�@,�ƺ����W܊��� �Ӌx�{w�����NᨄP)wL��t�}�\u��jPmue�%[6�v��bX}���К������"?��|R�)Vս�.�{�`:�*e�����eBƴ� ���X��lA�������)W��`���DM�i`(b���@&�1K�)j/A���m�P����j̟�Ŀ�}
��>�d_�h���Wp�Uw�'^Ey�.Җs�����ӧ#��$��e\{�x���pⱇᴏ ��rߥ���}�	,[�
FGG����1���~���zŨ�?��Qm%���q˽�#��&,��)qJ�ɪ����T&�Z.��I����}wŮ;o���g!�M�}`Q/��r!�|>/�uU�v�l6�l:��B���gL?��>�g���X���`&2��@:��U�,uK��Z!{�@Ӂ��j������ق��?���h��͌���nnH�#J̉��FDL��̋�Z��|��	�f��)��$�|G�nP�3��q������&RسrȚY�+P���V���>��	?g�Q�ijQ���`W�oH���+nu	����{��(8K���TV��o��5v��׊h"l�?;Y[[���ʽ������Qc���`�^S@�7Z��Q�y��:������f`�`��b��a��8
�:�^~S�*����W�y����Â��    IDAT�Ͻ�痽����14VE��F���>%3Bs=����ȌtS�"=��|����
$��������`��)V;��3���Qɵk�+��
!S�c�5���(���=�}}D�����̖ �c��}s��_0B��[��T��/Z��H�x�!0�%D���o�Ys1W݅��SJi��׮��sO��aP�+�^�LPw�S[ġ����ӨS��k�[LC�Fy#>�����Y9-�J�c,���(�'�܅7�6Q��Њe�Q�$$�ҽ`�^���R��bj2.�	[�*ֿ�
���2��;��,vں���wc(u�o����Л@~:�:�c�vr�^���Ɉ����h�fΘK��(��bh������,��&�5�v�udc1�:1$jM�G&�&($cʘ�s�XP`I�V9��5�� w�M$���8�Q%0-���Lb&IP0Ɣ ��4,�gKb$����;"�OΘfz{ddS��"�R{��ԓ�@f�\�n�is�,�)��1�_�)�W�u��K����?)I�Y�8�c��G�0����]�{<�ȳ@���g/��ٟ�n;������A��T�w��-w^�u X���_�׭x��eh���.��"3ҩ ����v�?8�dLa�~��xc5{H3�f�Hg�X8����݋i}�3i
Eժ[b�}�����8�}n=���aT�)��r�%/�Y�k�B �*�c�D�w���^nXmw ��|J6�����Q]'�Ǜ�������w���1���M������^	���x��ƂPPi�'eR&g�� i�Z^��w�i�=��9��3��K3ꑅ@���+��Ш�ݻ)�]א2&^F�`i����C�>�3���_��v�l5���a�������9��q˽���7!���l�ݮ�L�kd����a���kV��C͞gV�(,eŋ3iYyRMW�e����M'�(�`�#�f�.R?�6��%1@�:#zeS׏&.�U';oJ�[�*���!�؈��(|��=їnH��d7��\�_^v�l� ��a��>lZ��,���O=��c���͖���m���,����]u�=�n/����FHAz�#E��"(���#� �:�]G��,0��!�(��tz�@(�H��^���9�>��?~0��{��{����{�����=/bw-�2o@2)R1�,PV������I�����A~FZ�j2?�{;��W��b訋J��)�'��SeB�帘�ѕ�=�/e���f˘����.�8^.#C�i�?;Mw�C]�S��b#�6�3V�FB�^'���V)c|l7j��{^��8�~����xa�n|��ƽKV�<ِbg{ŒU{���η>���^T`��6�t�mx���q�٧�}gsV��p�����;�Z����	z{9c��bSض}���)�~<�F����&e��G*?���n��%aKe\���U����+�z����ۑ���5�YDU��A�U�!�w�q:��{8�� �岗����Ǟ��d��𮷜���=�Q�s�Z����z���@�6�L��ɾ(cj��3��XH�"�G+M�H�Q��ޣ�\�
�O�4�t2���i�
/.����'��\x/�'��ӯ}!�u'߈����W��ͫ�U�զX��K���L��{,�t�� @
0	hގ���q��0v��G�C�K$�a��c���if#~��m4 ��$�
3݋���5�M��������'�z_�5�©'�Z,�3E�L�Y�o���E4�Sh�&��R�2^3'N<�z�k0<Du�*�5�����(�L
UlJ?`�(����xv�<���x��5�� �T�=�H�{��u#��R�M��M�33�Pޫ�aO�@��r�E��y�]�n�Rs+a+��Iz,�b-ľ�0�������"�CD���X�|^�ӿ'
PCpf�`�^�3�L0��g���)�,>	0
�k|E<GL- @ġ(�-=2D��j�#,�������%�+ ը�����RoO� x拏T�{āi�.�tҭ�*�|�+�h,k��۫75�ߎg�L������N�8_Lb���JC-\�l����e�hV�غa=S;pʱqŧ/ā��U�M!
-�_�#�yl���hgtܥ�j���@���H)��PXE��͖�6�'X���cODi"9� ���pH�i������6s}�SH�����$E���lQ�q�Uiq���#-�'�j��S�<g��r`'Y�i;�Őp�R[�5���Z��q��REZ�=�HѕW@�����jj�*;(�&K����U�1�6F�1� Z����~��0��on�G��w�����-�;���Ǌ;'곫G�^��|�f���q�ϐ��̘t�r��#�]���&r�b.u^���k(ԁkox�{��(�2����&�)�
D"V�qG�~���My8��P"��|�7`-�DZLm�[͟Ӌ�ge1ԓ�n>�)e�RA�\�`L�����?0�|W��V�4�Ԛ�Hd����LA�{R	��L���s��I�%S���g� i� �4;�S	_��s�~*0%�PC�YD�5�/}�8�=���Aضc��>�
������L��z��z��6�A\$]A�B�
xb�� p����א�RS�H�XPuwV5d<1S��s�T~�-����&��&H���j5�:����n�vکHd(/�aՆ1���'��kQ($�gf����W�&[l��󈁮��e�t�Ne�j~I���YY��#7u��T����V��6.mWf��X6�g�
< �f2�7uLLlGi|#�~���ć�¢���T��_�\�_��n�Z�(Jb�59���n��-�������������W��Y�[\���*\4>2�#�x���d	u�RƑ��`/���tǦԓ�F{m�>J\Ș�KԦ
*�%������ 23�P�[��GM	�2����<Ӓ���MT�&�T+|r�Hu�������z4�D�_�;F��pV7�2�H��ݻ��R܆��c��~o<j�&�;z��M����e���$��X*��p� ���/�o>�$�yw[���<���s&�;�x���Xi����[o�K����fϞ%�d�r6m�M7ߊ��^���J��� �~f�Y��7���Ϯ��Uq��R�lR�4��ٟǛ^"����g����شq�Gw�լb��98���q٥���Aw�B%Y�q`�x���-xq�����ł�>1d`l�yt�.|�˿�ڭ��g	cJ{>{�D��2��g�>_��%�D@�@�ȸ�i�F��fhrF/�q�<��bM�Q�$ ������O*�����Lv�2G�^y�A'?bm�-�L�vŁL�|��q5մ��� o�q`��|��j8 �[n,gYs�v�Q�T��%	1��/eB�-
�f9�u�s�d����4N������S��:��=��c�����]�c�X���g���S��.T�w�?�Ƒ�SN8G�?�{6f���b7�6�F.�?A�]�����M��m�*�-����M<����}�����a��F2?�t�0�=��tqL͇4kWOu#&�AFJ�p]����~��(�nc��~ZvȔ���]Q`ʧ���}oG��[�^<
��V��Ȃ�2��5��_��5��B�|� ��z�6�)OϷ��E�a*
�n0&�In��T�fӕlF�F��-���*~6�K�7�AaØ����xʡ+#d��@���j��f��$P�{N;_��-��S��L���U��n��uE��9�3�}�16N�=G�B���iVh�;ݹ�SSعy3j��q�Q���O?r�y��p�|�����Jb@�JSe�_�Je1$��F����oS\Xđ�����h~DW^Jq�,���TF6iN�6�x��4UF- So���{oTjZ� X���I�T��_���rD���򖊘C�Q�n<�џϦ�J���c�Z�:� ���rU
X���$f�d��J�Yk�W��bF�+1hj����6T������0�d�u���"����sk��W��K�������y��Ȋ�%�̋��ͫ~�G~����o~o�����h�b�
c�)l����ȡ�������.ۂk~�g�zy��Ӝ����1}�|���?���.r�˷�+W݈�&��&���ݝ��G�sO{-��?�lظ	���׭���8*���P~���8���0���`g��>��Fj@�G�E6�A���h�NX��� J
����Dd��TVv����>�o*1d"ͅܒd��("�2��%\����{�%LnX�b~��k�{tJ'��|�?�A�ATMy�a�'3Lb�p{׏O����G�y0��F�J=�$Â���3���_	�n�2��a#�m��H���?mԯs&��(��Y��'>��O:<�ŗZ�����n��/����E=F��S8���ZObl��O��S�M��.�{����6]w9~���?���z��*�2�Z����4�GF�DM�|ظ-V5������v�Z���73�s�x�<p�����K��u#���151���1	*��6c��<N:� \���a�LM�jq`�.�oK�ۆ�������li=�Qt �(�`�l#k�i3�DCd4���tBP�}��"��7�,�P�*�-�_:��#��-���x[�����e��$n����$�S%��r~��K�8���Ҫ3�'b�"�J]�Rq4��l���#;Q.lì������S��b��w߱;w�������c�9���7(1lî���.�w	.z�98��G�<6��yv��<�=R��C�lꚵp��;�f�z,X��pz��d���w.�?�}X�F7�Tj$RL�x̵ЗO��}�ĥ} ������^x�E<���TJ�o�E8�=ga��C����u�� ��ow���1s�9�X8�-��^����W��z���B�Ir&%�>M�4N�0�SO%�rϒ!OJ5�x�
3N�-�\��L�]�q4
���yx|�I���Ƅ���-��:-$��lnc$A�Dߓa��9� �_Y*�������J�2�� E�i#�� xGK�:�2��ݗ@��n��o5��[�d Ƌ^p�%���y�	����L�:���uh@3�<�6����� yw&�#0u(�d���M��M���AƸ�jhL�F�Y@w��C���K?x6�g��h3�N��<y�X־]��7�q�wp,��vz��	�(Ϛ
R��B��?�t'V�A�ՇV��L��]�r��4-���"�i����h�����ㅒ�	]e������*+�p܃�s��ӰZ����>�9�a[TT��{��a�)|��OQf����$����#��Z	�ǗT��(�סi���b��3k��O��%��1 ��&l��~� �GZ�9� �����������.�W�m�c$e4+H�'p�[����ES��\�k�4�����W��떵I'Z�}2Œg,J(z�@�P)�U��N��c|�N��؆��w�|�������K0�cY>!��g��<��j���I�'��PI���H��- ��>��E�o:^�Æ��,��	��J �ۋdO�0��59/t��94?ʰ?��2)oY���g(���#�M)/Ku��X RZ%�ȼf�E�RIr8�E1'��*�4��S1>
�;0�جz��	Q���c�>�Ӄd6+��b����o����d�+��X�j�����1ݷ_zL�S�����驫5Vo��4�X������������1���l���c�mRާ_؉���xp�Cx�A�˫��s�A�,�E��+1R]�
�'�Z��a*%�k6���	�=�
�X�\,��(Gl�Gq���?�:V�8�G�ځ�^��Z?!��ba}�9���c���ށ�3�]-��gV����c���7�h����r Rh�����/o\�;^%2������b�@@�*����){�⮯*909��x��jg��S�����ixX��1�f=�X�X�~�O`��`�+�>��Z����b��q���Fa�"���v�_�b�
�W������J;��H�x�R�p�ZuڤnQ��H���$4v����6��EP�4�'S���?����ec��p��ͤ����,�9j?3��b��1�g�-ƒG7��̣�H�'�T����}�s��[�A*�h6���~t�����8���(�%%�c��.j�"�HK�TX�+E�2qwD$�h��u� I��^Ǒ1�
��"R�&��9�Y�]��(n#�a�4��7H�����^|a��Itg�8��Cqء{��;�b3�%O�Ŋ���\���퓊 A&͏�c���h��L[-�����S�T��h��.��q�y�6Ǵ],�+o�ř��[�����D��J�lz:0�h�r�q��zs��=�R�ޮ�J.�2�^l�g�״u/�c#(�va�@��L������@ 7�N�oS��cz�)�k��mO�������.�� S������g�]���(�x��X��z�ϾX�pj�֮ۄG{
;F����Ss!�U8B*Nd�Md�~�~8`���?ЋvB��رs76n܀�;���?��q�*�L26�?/~ +Vm�p7>z�P^�^X������;�ٯ�v���F����H?�$Liͥ�M���\U�F�BӢ���\��=j/�rsZ���� ij�[r~E(,����Y�8��d,�_���W����;k$�E.�\����)�����
@�M�y!��NKN�R\Y0ϑ�Cb��%;��{��BvN��C� ȹ�"MXH��[��~f�=u�3�Vq�g�MrC�737Ŏau7>3�>�~�y8/\�,�v� #�fv�r�"�����c��_�	k�w���N��k��nYSΞ
i_�2�b�X�� c
e�dn���<���	<���Y��D����A.-��=�|k��4O[s�y_k��dޞ������wcQ%Y5�}����}�9PL��K��{~=u0w���7Ջ5q"ҿ�k]��+뉷�Qgբ 5�\��� #�k����j�B��i������jT*�1��	���06�:60ᔵi�t:H���V�0��]ܞ�1G!c�hVЮO!Q��o<W\�Vgu:����+��g���jT�#���n:v(� �:2Q6�2�2�� M���Q�C����'�}��q�k�I��='����߿x=[9�vv&j$��w-9��j� U�j�=��)�+[A�c�'���m���n�6��y���I7[�ʛ�X��)�'����~�q1��8�ƳI��1�RHb!��;��f�b~T+�D�+��ܿ��9Ļ2h&t���)���Ϝ����9_D�VU{�	L}ޫ+��!�r¢�/�TS�jy
3?:~�~|��
0��9_N�'0}rm	?�����rL��3ԋ�>x�=�8W����M������c���?
?�Η0�������/�\�z�[�U�L�6��d��F��_��n\��У�<��Ջh5'�1��g1ԣ`����gv����Vo�@��2�qu�̷�/^���������zIzX�)��v��o,���I�m�*��9���"]�e3"%[ڤkh��z�&��L���UM�]gUJqJ����L�@c�=6)7*���+H�9*���l��Ϗ��s�Z�2��㎥��O7�\i�A�Ä@��o?`��-`L?o�-O�=�9��N��Б�Yr%��V�9���E�c���?l�@z@��H������m�ނ�fI��d6^0�A�Kq\P]t�� �ȇ����N܊;K���O���j�Z]h��z�F<�9��WQ4gm�˜�wi��D2���BS�d:��ܪU��\YtKN!C�/�x����)��E�a*�� �3*#��0e�|聮}(Z)��O�l4�S�~Ε���<4��
b�bH!�̨+a�!@������o�,#�����3X��\��+���5=k����� S���d%�u4�%�X�+�=�9���нX�^wl��I,����e    IDAT�Vjh+L�"������E�/�V:��IAi�Ai+��d��R^Z��L%�[���-� ��r
����]�,ѭ�E�-#�Z�"�=��1��֣q�{��U�%�����E�����:�{��-]���]�3�t��E�
��Xڊ�Qk`|�UR5����C�.~�ES�����)���M�#]*54*Eq����jaͽ�u�&'���S˱���a��Yr�xэ��cǶ��[�~O�\���<.;�T�5�U���r�����n��B��������(��oP��-�䱑`���&%�H�-�_�pjl�$��6
�r"P�k\zg|?N?L���������rCB,�g�E�"�������3��ā�Me"ū T������QF��S�&btaq]*�:�"PD��$`*�}K��q`�q�c>�=a_|8K7�Y��uj,���љ���K������Pu���Ռ�r7XI�M	��M�U�v��g�����/�F�.��¡8.~�[��żYʎ2�p��w�E�gl?��1HN��cS(��C���^w>+��3���� '@ؿ�/kE	q�V��gB��~������x�~�3�]`5��|7����'��nʀ1Ig�����|��������p/"�v�9���y��瘞]z����;0��r�^�Q���c����>����^�<l�Lb����.�ő�����-jlV[�ߜxp6-Ds:�1z�+'��+M�k���b��a�Aj�z��(�YV�����,r�̰M��@[��{$Gԏ�kLsY5��<J݊��1H�:*������Տ�3�cjϗy�T��*����r?&+�ԍ:�o)�S,Nj/��o��s����i��hՋ���	|��7�S}?��H�D�g�O6����z,_5�fz��$R2mA�09�@	d-�E�X��h�(h��Ѡ�A��0���uNĠ���ˀ��Od�Q����iB0e�>��G��K��<(_���}'#���S�;4@bN�(�Q.��H�	1P�#�ϊ����|�gs�g��*.�GdL	L[��|=�ݍL>/`���K�8�dzs$�>�@�T��������q���q��?cZ3���5E��ڛ��g���=����w�q�K0]��*\y�uxi�J\�����^����U�PJ����`��+�ڂ��ҥp�����	�v�$FD����y�<\��Oc��Iy[�_���X�~5�ǔ�0{V7�;�d|��o �ErgG�/aܱ�����J,�-e�7�.Ǎw��H1�l�Get��T�]'�V�4P���zS�A�oj2��A@
�NA��C�@�
B�&JTn6sPx���I$ۓx��C�B>��f��Mx��g�q�f$��c��Ő��t���P�<ë���R+ϩ���5��l�:d�^^Z����݈�+��X�&av!k�pg�)O"o��ώ�pS������v�bk�^P&�2�8����7����Ì���{�n;�_��5{z3��Y��zKe9&+y:�K]�T�A��5�ˢ�[%�d�ɔ6XĠL��(�)/?!e�\��ç͑��ru��9�B�3�"
�5�@i����I�R3*�1�P�J�le�(�z�fKuqf!Df�e��!E{�f�<�4x�k��`�
<�j3�Z��XFe��R�˾\�:Z%�1��TS=4?�iI�N�6�Ձ)�x���V�Ǵސd����`/�]��8�YYɚ9�5M�"�T��4DʋR)�Z#[Hc.q�ӞY�^J��'�� ���tȓ��v�'��*�XG:U�{��3��k��`������_���k~s3�-[��X_��8����Z� c$�ҤN���s���;{�,陏���Be~y�"�d�)e�ڼwU����"0U�9H%ӭ}�}Ke]�|�IR�f<��&�z<�m��,ǲg�`Fo=��X4��Q\�T�|b>s�o�qg������\�3ۂd��(mJ�`
 �^��䊂if�B��-D�O���OD��A��-%XZ���V41u$v&�s�����v�6��f�x;�M���{V�}cL�.���T�n=eѱ0���g�="?t`�ܙ&�z����-.�
¯#��H�O��1�?�<���/���	�Qci���2^�{ʇe=ʦp��,ݠ� Q� �ejZ�cX���h�^D������#���F۱��& o���ʤ�L���7�`��g�r�:l�5�b�
�J�_K��4�/u�P?�>�`��ڣ�h�0z��-��E��Fy5����V������~{Ýxi��3� ��h��$��s�Ga5�tQ'����pƣ-l�����y�'�։�cL�5gL��R_^�,�cU�p�s{X aD�����`�� w1��A$\WA�OcE�P8�F����`S���׸��<�QIx�L�H�������rB驂)_�G�T��J��M��"#�����B<;����~Ζ*��@�yU�QE�:�Fq^�k��/���]PGV1zb�$��V�Ǜ��3+7�X��*�z�ZM�Y�9 h	LE�C���͜8����'��>��t�3�_\��|b�+	���/\��_.��B�y���������F�L����r�X}�����16�0��A�+/��¢Z�Ii��9��J��j�Ei��c&���]y�)�Dױ�.d]ɘ����\�X�g@��G�i�>�0�"{B�i�VGc�}�E5x�1gO����4I~���P���~1A��8�,����E$k����=��	Oh]��j�ݦ���Lz�y�3�轧㼷��9���������a��5��e���.:[�Oe�۠�0<�B�n��=d�4X��)�ƾl�>��c��S�=)c�p��s�>%,(�2�ÃO�2W�I�kMTJ�3��}�)��Eo����E�C&�E��S&D���n.?��c���0Q��o�tݽ]�K�9.h.(��Pz��}m�o�I�Oתo�(��K�Q�xj�M�v�<�t��l���Ci�2�&�P��p\���QVd��X=ァ,"�T@�L�|�g�	�t�X�\��+d��!�����ˡI���S��LPF]K��ڹ^4 �;�#�W�_�@,=aL�d�7�[�F�L
==yϚ����ox�zq^��f7��G3Φ���|��2��� ���d�ٌHa	F��*�����5�:���v-^��<1b��_VT���9�b��7p�]��v0��@�6��YoȈ�J��bqJ��K�hӖ����b_�V�P�F���m\���p�oA�7tw�����i�JL��(q�6��i�L�E�&�P/*0M��I�h+��Fj�bR�`ZG�PAe��
ZE���i�Ó3*o��ׁ����ő�snHph�0�e�8���;� t�;�S����@kR$cz	�cxƐȯ	~�~��K�:��&˻P����s����N�k[��4tvfD�dM�׀8j�����.�M�/�����ov7�����y�}��l��*�
-��&�X�t)�̞�#�:R啲�� ���i�06<ܕ���e^�f�^+N�a���F,�	��¾4�x��Gp�M7�ͧ�o=��R=��[�ű�J��)<���dq	ӡ��EL�<����o�iWف����R��8�>l�HK�d,��x\��x%`��ch��ɔE;�Џ�I�<�S�cB�p[���ʹ��ȗ�<���Y�\^�f�Fc�=�HOlX���c[T���PL��X��� ��'�_�1W����[c�^?�:�j;�Gi�&"�� ��g{K��%r=�2e�Bj��T�h�>i��%L_^�в�"`�ٵ���uo����?a4_k6erg���E��x����;�EF�:��>��b��~����eG	O?�
�W��V���E9�P|�z��9����t9��6ݽ��f��k�8��p�a`ў30< %dy)�*�%���m�<�L���?�Ȋ��&���f�]\�$����X4l>�����ޚl����sd,LHTt����+먳��<hbҡ`���6`��'xf�
r6�~�,K�.���*-0Ό��H��DbO2ª�y�J�i�
N;���Pg_]��#�g�m��0�������=��>���f���Y`��K���Gaa,�ΰ�)y���iL�ͽa�6�5�J�פe�ZG�6���d���7�7'���Ә46�����q`���nW�	!Eh�5��h.*�R�leA��ψD5�h��7�93{�̥!�DST� ����K?�� �=S�NSٜ2�$)�5�+m���Qo�r���G�4xXq��R�K���^�����&��/��M�G�\C���sD�$S:ǔξ�� �)&����l 7K�s�+U�
S�H�ES�s.N1����뚠���[�8�B",�.�� '�c�s�8n����#Jy��X�v���R��ߠHy�SW�D�Y������O��x�9Ke̛Ջ��w:�}�q�M���<�?���xy�j|�#��������D�VGv�\f��jK�9 ,Q�C���W�q���v2���i<^�!�����0e����/_�G��T@��R�fw�3N�%瞂9��nش[��@�Z��Tmԑ̤0{�l�tw#ݝ����o�� ?�"��,24H����	0%�ʧP�6РK/�	������}L���U�'#A�e-it�IX1�YG�D(4�c�$KX�g?z�t�0{c(Mp��R��F�D�$2��Z���۫ir�vHW"��ƾ(�]¾�}qz�f`F"�he�$����ε���B�z���Daڒ� ��|���:��]>S���*UG���t�2Gh$��dKwc��@��A<7�v���h's2��O��;V��ٌ�u���Y4�I�:ak��
��UV'K������V16�X��ɪ�5Z�T����0|�I 8�O:���>]�9ʠZ�B�^�P_�fI�J�\���IS��cjb��QTJ#X�p����q���E�ƾ��6p��/��w>������E2�Uy	�=��v���2�}��	0%��G�h`�Q/d��1��*�/�Ԥbפ�t���^��TGfЀ)�o"�f2�	���b�2�<�J,l�?�0������@��No_����(�5��I��hb�R�Xy��$�"f��a���g�lteU��=`US2!�B�r�v�j�Vl�@�]ǡ�z�O_���e�Z?\聸M�2۷���/Ʊ��<@�ɢ�[�00�	{Ђ��h�:9&�#�ۏX&k�C�4��u׽��u���G�O��Hg��00��}O�g�
cz�٧`�P> ����yh>���b�n 78���G�J��(�UTk}����G'u�-n�Ir�;0#��h� ������;=�sws}��A�i�_ӏݰGU>����=dO��6W\���#Ώ�g�Kzf-�}g����Pֶ��"���`4X�'�©9�"�Uѡ�x \�L���*�M����[x�]����~��B��w/6;��bB�W(0U�7d�t �7q��Y�S؈K*
�J��qX���d	o?�`|���b�L:�S��� mZbV;G����Һ-x����䊗��]hǳh�)��C(�E��e��'��r�+��8��Q+3;�@w
�� 'w(N9�p̟�‫¬%�&�A}�&~s�]����hf�0و��W{���5Sg �����:b:�=�r�ў� �X��vh��X.������8���Yp��&Tҭ�Y�rY��i�UA���P��>�gnK��Ǧ`�����^��s�h}�s.�^N�ưϠ���kI�lmP���_�=��L���] Y5��{׈��t+H�̘�F�D�m��Q���(�zSE\r����ٯ� M���2��?�b7��k!)��txfj-_�>rU�W�3�8������
p���⺿܋�JZ\��-�E�XB��MbS�Y��b�|?���-�9�f�����V:%�G�|NS�ᕱ�k:����c��4e\L�m7u��m�e�K	��d��� p�E�TG��x��dL��a�bȸ� ��A5`�M���˙�<�(%y&&���x�'������Sk�%.SJ����K2�R^J�I�4�R�[@�6�������z� �.{i?&0}�Y����.~��8紣їU#�e+6�G?��W���/|>|�T`I/����p�ma�*�BP�e�+����)��k˸���`��:b�� �F�HU� �}ӯU��܁+�w�l$uL TGow������їc�R[�nǃ�>�����R)#���X�"��`���h�`���yw	<���N��N�Κ.`��t	VD�k���	�Sw��I�OI�0<��X�M�5n6��F����V�x��8z2U�w�)X4oP���X�,V>�"&'J"�S�X&�J��{E��ȓ��D���� �k`�!Z�9 <xG^�'�ae<|O��$g:`�`+�6ʔ��x&$|]�@x�ʷ�h��y��G��hUE���׃�
k�L�Qm�0Zl�M�X�e��0Z��i�D:���.�w�H1��lKnr��J����5=��IA�1�v (�52s0�G:n�Y#521`�,�8�ف��r��Ш�P+��}g���9}��,�(8f���f���R��05!`vx��{ �������Q �.]��?���1�Z1�Y���M�k4��lh~D`Z��ǁi;���������90e�#�[�
cJUB��B#�q3����:^z�i�f=��0��V\��6Œ eo����n}b ��<d<~)[Je��L.�L: y��d*%���R�X�Zh�A�G�UB�]E�V����L(�?X*�T2dQm$�(�FO���g���\��f�䠐����6�ț�M�a�&,���x�N��E��oӡ�j����:r�<R�ãp���2ð^A�=�-Jl���1�V[�8�Zw�u~��?`�ޯ�}��H�|�
P�ű��~�
<��˘ћ��u)(�d��+0�2eL�ĜA���X�U�XD@y��
�=;/�I,��!�OM�צ�z�����	���Hb�,M���!)��{#"��Y�H�桎�h�x�R9��c|fK�C�T�-�{�j���0T�x�ѕ��I2�J)B�ǏB�h��y�Uǅ�����E�H���4������k�xo9{Pt49�0_����AFn>�㡣��xϕ���Z%�.�����̮&����p��âa��&h�A������� �=�?�+Wo��]��6i��3�x<-�R,!ĳ��8C���yZ< �P�-b$�=���f]��;b?����p���b�b�R��I����y֚-m��և���V`��C<7�j�-	�E�e�\�]�tO��ц� n�RM��)�(�
��>�̼a?���8 ��� �vu �8MK�h��=�a�ѣi��|-`��,^��bGGa9py��e3l����Q0i�"g-='�1�rp��C��e�[����8*-+�:�ԑW����Բ7����.�fRm�6J�q9����{v_���8�Ȓ��p��ӾN[/�z*��6vSe* Օ|��/�O $?�1������+�p��܂��Jh�zьq�|N���:RP_)0��&'��#�;uH*쀐�=Z���tK`ڕC#��T�Vp��
L�tC]yi~D`JEV���LqaL��!mO<�MN��HR�3`*R�2ʅ����x=^�\Z]yť��b�M"c	��C�_&(�-�]�J>��"�Bu�yJC��kZ!����;-T+�1���8���Z�u�LY�~��q�1}�Y��U�5�\�N���#�k������?��=����.|����9%8J�2`�A�+N�՞���ƛ��y�@�_S��>��a��J��l��nM��C�⚫>-�)){�%�m`��sL�id���C]�?܅x�"}~c�ؾk��AL�e:RIt����=��9V�X��dπ0d�h"�̕�����&0�!�E4"���h��*~>��]e�2eAɫ�����p�&wl��Mzl�ȤZ�7'�h�.|�+�`�W]�(M޵{7�r�.]&:}?P��(�����T%�pY�U.5�i��*���7aŽ�'Q̂�UK�#g�    IDAT*�-���D�>F��h%�����7�n��Qbu�T���[-6�3@Ӷ��x����:g���X�`� ��rX���?��A,{i7���7���r3&k���ܵ�z�r�bA�����Y��`'���\�LĞE�A��d��D�cK��V9���T�>�}'/ь�TC���=�D|��b d�1��@��<�bJ/��w? �bL�|�K����c{9�bH�T���Ɗ�Ë%T�1U�'��@���VY��@+�!.�7ъ!K��&��4Obc>6��� 3أ=��ʫ3L8��X�&SH,W��N V*	�S"cKy�	p����L��3�/ݸe�	GD�\�#��|&"��R��\Y�`?]�zI�tI�P��k�����d*�X<ĕ]O������w>s	�Nȡ�������f#��׿���_�c_{��=*0e�lr��j�����l�\��])�$�WJ�����iH���߶�F�\��o����zx�A���[��������<�eO��`o�u[l�G�<���ʵ�:J�{��64�G&xϯ2.����	��2�<D���z&E�<��E�O�d���?��Y��(���u�_��J���
��aڢ�%�Q�y,1�~F�5RY�'iѸ��b"㎄1�B���&���U>�"~��3P;�`����4�S�mQ�4W�M��%��e6�jz�I��U!{��R��٦= ����Q�Y�e���Q/~ʙ�q���W��zy]�)|�]'��3��^ ��h��G�p�����[��CO���R�D�l7��'}�,:%Ua#	5�?�B�ມc�A���,pIN�q��j��fe
��$����w��}*f���W��$�
I����W��-}S�.4�]b
�EB�U ����Y��G�%�f}O�#�?M<��%� ,�ߝDE�����d�*!舎��37&R��z�3Y�< j[�H_��.��s���w;�*w�2�*~.$&j�
_fR\����6�|���`�Opo��`����+���8��|�XD��e#�¼�
�N���,ַ9���v]�1�p�|�C���{�@����`�BD�!�i�༛߂>j뛵*�b(5�'W��W��>�t#�'p�~������t����8��_,��>���s`�~n\	Lcy�|?�V��*E��C�-�G�Ru��+�P�*c��jW�94Ro�3�ա_��h��d^��;6*QP�-WG?��<b�ZL-���S��i1ך*�U*#O�h:�I�H~%�2� ���`*cgU:����h~�)��\����>��~z��x���T��{�,aL�z���(�{~�\yͯ���p�i���W|]�;��[}�<d���E6���r	V\�fL.���{d���k12�(�}��*�:`�\���1��ߌo��F��ɀi&��X��ZU:N&��0�r�c���m�|����C��Ď����̡�ȣ��"��B"��h����\(�l�\���Z��Z�<J�*�v�~h�c	�%!^{�ʊ�Ø����CBd�%�5'����Q�j�q��w-��~*n:M(��'�\~Qe��C%XPA�7��9N�p`[�QPvg��2O�dcvH�#�e������ 8���V���z�dEzfX�fE�!�d����>�}�;ݯ!8�`؟�d�n���Obw9�j,�22R����㢤�fXti.�ʨ��4hd��d��"7�����󱊝|�JF�hʞi���MЃ�|�@Y��H��u���D���]p*.~�q�2�v��e��������T�{	���n �o5���9��v\�s2٬�XS2�h�]��42���v�^��\JS�.wS �MPG�u���T��%-赙?�׍��um&��b�l�����i:��k�����������q�)ѕTW��e�V���V3�$*�
����J%�+%:���� ���z[*��f�JA>.��̸{!���)55j@����8��{��{πZ*�����X��m�m�;^{ܱ8��#���5�h`jtL��|�˪�	yF��lFr�ZFal�T
��ad�D#%k�C�R��n�'�����G�������6�H`�,��y,{z-{r���'a�P&��;X���:lO"�?]�3�da�\����@U��4o�J]�]��,N�:#��&��~-QP�@ȓ.OX��D
<�dڊ@�N`�.��ڃR��9rG�����CQ��A2�#:�g�[,�ua�y:����tϋ����&8�D)��Ҫ1����쾿�3��6[�P��z�q�\�-��;4'B�D�*���[PlЪ��
�H�S�\��M����d�8˷Q؁#��ŷ?�!� ��4k-Ы։� ->�W���X�u
��2h�0/Ev�G��0f&z@�A���E`*��u��ې{�w�D�ZG���X���h|�3p��>��{jL�.bm4�s��������g�Z4�3�"8eђ�0߃�����o�l���\l�~�d���:�i�2�V���E5����Ln�A��(��y�^�gG��k������Z-��3��kg�}�`�E�vhy}�1�S��
��F@�ǀ�{��H��gj���^$k�9h-Y������H=���<��#�d��܌���.��fL�bI�^E�-.�	d1��N8���=7���a�[!=R�Ҝ#{�D���mj�A�BS%�h���e���;p�c��J��Rټ�,�Y*��8
���0d�}h�����{D�{�jG%j��P��G���P�$y�d;9��#qS�D]�i�A@B,��-�kS&8c��m���r\L�ZE��U�%ө����	ɹ�{*3U��D5�0���
4E��e�o�SH��O�y�}�{k���m�F%2n��ժ|�%��8a�\q�^1.&���zL��}i?��<���2�t�����ޤ�)�kw�W�ܿ'q ~��oc����L� ���o<����A5��P~��~wJ5��e��u�c|�0�����~���-%I��^�tgo��*�`�?�ysfb���He�X��F<��r$�1�{�ix�i���7��
�z~#n����ZF=�DI�Ɋf(��fh_�|�lV�z3Y���+��#�C�����QE�ȁ<����Y9.[�
b��i|����	��e�R�߇�r;*��L�!��y��6�NB��ڰ������^�'�����#�at��=3��=�"	� ����q(EX�>9�,���T��'�yK*�n"�h�������F�� ��7�gź
���3X?�F��D,��
�X�K0��)sm�:T>��$O�lN\zɾ��P,��T��\39VY7�Z�~�({>}~dau���}v�]%��֛42���V\~ћpѹ'��*��u�y"����`U�a��SH`z㽫�1�UͣB�s�ÖC� �C��G�Ѯ踘\?����KR��b��'���D��z�ɲ{�^�؜�HH��S�d6{��hrϤhJŀM�NS��qĊ�K����Ss����Lɶ��TJ���R�qZ��J�6q�#��*�F���:�Yf������3Lti��Jd�U�F�v���l�/|�8���/���B�غq;n��8���qđ�"AS�����Z�Eq������t�V領m�p�9��C<�B��R�W_i#H�Rn�[��_��W8��c���W`�^�z,�q��V�'_��@7.z�I�g�����X�����>�Bvp��uhxd��m�'�Ar(E;-������0�:/��W}��*9&��%'��=���H���~�Xi�����],�jQ镁L�?`%rޛ;$;+�X7"���}���Z�7��[ �Z��t��Ք�$�P�.�@3��x�f�P?���*�@xP\�!��k�6�]���\3|w늋�R��~�
�B�-4x��� ~FR�"IP�1@c�)LX�e�T�|��8��}��Ϟ�9t��SuQl�cҿ�m���e���'��
�1&�]���d5�U�'�@�^J��5Z�#��hZT��.CV �y��M������ʻ��c�Ň�?��=l�¥�hm�� :��������U[�h��?O
w���������%h.�W�βK'����ƈ2������3�H�b��J���x����g�|�?��e_���kk�N���y�� ��[U3�k��t�~5)�݁<d�_�Y����	�9_��h�aF�Ŭ���-����7��y4V	��1��'a��6�V��jN�1f8紓���ތyCd��%��-�k�+���pFé�U<"j��w���.���UZew!���^1�3�!Tt/i�Q㛞2T�2+�٤1�L`�3M16Ѧ���R޼�r�Tς��1��s�r��)T'���#xTW�nĥ�4&3�%?4��2��9e._��	*�����tcʞՆ�y�+�3l�b��RIS�+H#�|6�t�dLU�2�$Y���	J�s�}�2��Ҫ�v��t}�"R�p��|��i�>LWM�~�W,}�)�E�f�L|��3�7 ӗ���\�%K�>s��+��#��8�`�z��+aQ���}���r+�9���4���q嵸ﱵ(�ٯ��
9�u
�4?���E��je����|�꛰~s��]�$2�2�ٳ���r�k�Փ�<��*�x�b}�ax�;N�x0oo� <��������4��bk�̦�5�\(`ʘ���Hg9)4�aoe�X��I5u��f�O�k��kA��X�N$hxP@2QC&Vp��O��5#I16R�?�y7��~T�ӨHF-�m^�J��7��4E2�  E7m(ٙ^�����0�w$.A`A{��s/P��{��n��z�y�\֘��{n6P�U�1m�kx�9��y睅|�t���(C���:~����y"�v�a�u�T�\RU��Q��Uk��j�ϣ����}�2r��H�--W+�l&�%��Fh���H�<�\y0$S�&�ʳ�+�����&v�lE���~���>�6�$d�Lyn�,�9�-9����6����|����奟*m�)�!G�0P���4��Ǵ%�G��>aL�4R���1�a�I`�����RE�?JIȘ����Y
`0eE����/�����j��O0��W���0`j�\�T�m܀)S�&د)&F:Hz#�1�Sϰ*�L�����e�(���(�J�H3ENǂ��K�ᬔ�h�����-|��a�^��.�T|#������1��o[�E������4�r�Ԧe�[I�l�#T��V���R��L�*�$�ñHI|�
�n�y1���:�z���?�#i�(��W�	0���+���/`�P/.<�$�9�u\-t0]���ʯ�m<��О���~^�,6Y��˸B��� �DQ\Z��G�T	c�飻��:�LT"�P�z$/�{f�#\F�y��2IѨ*�L/E ]�#��L���Y��2V~rD�y��N6��p�g��%`.���ׁt�V���֯L����MK��nl_���0f�9&h��a<s�r�uz��=A/����V��p?����Y�~쇸&�u��И܄sO= ��ܻ1�\M��!\��Ɓ_��^�v�r�.�ьw���nJ焲��9�g���/Ҋt;(�kh��z�9����T��˼���.Ԧv!U�a{�ƿ�=x�	� �P@-m,B^'P�����ş?�zr���`|Ӣ���%E�ޫ�<v`P�6�7�Y��<����Ip��ή�v���{ξ1b^�5�0'���j�L~m�r3`��&���H��2-w�s�
Q�/��=s�r�0gvńn]#��[���;��\�]��(���~I*��k��%���ÆuZ�=�EVݖJ�(����=�lI%b�U�P�LH�J�^B_����r"N>�pt�НI���s+T8��rQ�������������x�
��
���
����s�${Kf�����NK2q�?��ѭ2F�UrRq��J�z>1��Z�$.z=L�d.S)dz9+8/R^)V�1���g��� ���$j̓Xd�M���n1?����>L����:�f̕��)�Sb~�k'�tWΜ}�R<�^�P�~|�	�6���QـiVg��Y��۳\
���N�]P�Bb��D��i�F`:�ٯ߀iN
���ܱ~�/2.����.�~�W,y��0}g L��Wm�U�\���]��t���%��{OG8�yZODr9�I���.�<���r$�|��Ώ~�gV���.d�2� �)~0��a�%���w+�}�_�a3�.r�6d��C|����"�S7щ��/c��g�����=�!��2z�}$1`�3��ތ_��n��i�B�֤�\p1��MmC��Hft,����GLE�oʹ�Iԩ�v�h�t�����H��u!��d#i��3�Z%���k�~�8�P]�(`��m�ߘL�X���X��ρ���C �	��($D�\�^ō�W���hEqz�������w:p~��<�KX�&
L�����Ѡ�K��y{��y�G}$M��QIc`�/���Wb��G=��%��N隐��J%%�2u(4�1��l.���~�]��*UK%�%�֪��)&�s}E�S�*Y���@>CZ��34�Р��o`dt+ڕ����������g7F�nեJE�kǑɦ05Q M 5s��}l�W�/Cގ�����%k���G�GcJ��9����^�.�������g �߃F.���D�����9�i��a��Q�(��9��aʡ�8r����*0�$���L9ut�rUz^y�d̏�E�1�N�m����P�21�Ԫ(V�0��艛b�y�c9d��-9B����X�-6.ʆ�+b��&b�:R�*�c�o��]�!���dL-�^);T�q�K,]�ĚSO=�,WBMG�H�`�q��	�)����_�g��L���a�Ӄ�Nj�կ��;���_q�Y�V�ӈ�0Zs`�{�����u� �w.]��|�����`���2^� �Y�B������� k�}�����Y�bDQ�;�rZ�mb���`ƫ(V�ǜd%�^��zA֮�Pkg�Q�x"���Ϲ����3�q�d�b0�~y�Z4�
RU���}u�^�W������1�AA���?�����[�4�[���]F��8�"�Uz�����,��L����
�$��(d�u���f!RG��e�`��Q���(��8��a|�sb��j'��8�s��տ�=��A3=�f�9��(�O	��}*0��֧&�PB҄�2*aY~7�	���y����;��T����n4��@y7�����^���z��hI��8��D
۪��W�z�V/�q����8���궧��U։���)8�mIEs��H����CA^��t���I�����b����N~�:0� ;Q���93�s�N��^eDz�-E��Y�280Rɚ�c�����L��8�:�ZgN�	ȃo�kvC0zoȌrc�u�xCs�����pJ������-ca����>��	�÷8X����j#@i�R�2rɘ�I�e댓$��L�sZ�O�|]�O�t12u�-�j�趱�2��Ħ]��Mv�&N���Vw����km<b"����ika�V!l�Ѣ�G�/l�ӂP��b�u�r�4'�a�SQl��S�J_�RM歓ؐ������.aLi~D�"�eN��֤6��'�4�U��Li��<*��@)�;OY8�~ �~!!�9��:�S
L�zY2�����HL��h�� W��$(i���z����O��ˉ|9b�ֱ���ה��oƽK��T*������|��2���t��1|���a�Gd���������e�c(�3�"r���23�����+
��4>���/�_܂��jhź�LP~�*L���<t�\�� ���"0��ߌ[���A�0�\����_��8��>y'�ε;�xp�S�����A7+�V�;caWm~����s;1U��W	������bs�    IDAT�Ugy�r�������fK�D�&H�bEX�j�"A��3+)�F��O���	�)?�s#Ud&P6�D�7&ЬЬW�E�HY�%S�d��Y��X��2+�H���#hZ�utո�͟hX�s����܀�$K�7x��qY�?���ϼ�7V�zP�� ��e&d:!R^&�jIu���̙�}��s�����RY�ilo��g6`�T�\���cE�=��=v`�Yt4��c�Pd�)�@w�)9��&'�Pa��9�I�7'I���
�N�b��FW]�qE�'~d�(�ۆFq3.>�D\����������l؍[o�����S��`��x��`����q�Egb�*&b	`[������Mkv��&�QPa��)��B��)q�%�Bz��4�g��L(�_��	L�2t���D�����8�����R��4�T�W��Lkc
L�9P��#)).i�+�I�����K$��S:59`�fGPJ��2_xUQ��`3˒�a����W�!ެ˨���8��㚯~�rӁi��K&T A&�a�Vlټ�~(�z���f_� +@Կ_��M��J)�tعȖ�R(B�rरm�(~��넅��'.AoWV�4V�YE�%d�����e+Va��>\p�	�7HC0��R�B`�_�v���\�0��dA�?�����MU�wc׭��>�!F)dW%w����:2��`���H�?��<�L�X*��2"*�[f��Q�j�Tv���Q}�Ng£?$��HcR�$�({�a����,q0'R���?�y�+UN��$�w0U���T���������Ɔ�7���1��2�5ʘjƠE99}�ET
mRE�?vG|}C���9:*�h�hA�����R��Xm{�6q���',B7=8j���E���p�cϣ�E9$R�{�^n:u6�@�)�]c��ڌqscuj2��ڽ�ǑQ�)ؑj�Af���?d�UZlY��^Cub+����������h1�[}�RޭE��7,��x���� �����W�tc���	Mj@A
*(~���pt���8Ψ3�c`L�@�Q@A%� �0$44M��*�9���眪���}Z��nթs�w�{��ڽ�2d8�ы�!�=���U0���T��D
��Ai��rz5*s�]���m�����D��Z�~o*cf�~{3dJ��OT<�O1���X�)��¹������g�k���Om�Dik���"��Y9[\��c�`�)V@��]d����q� :�+U��[m�+�D�g�(��$]0��3�U_������<�ۋ4��5є�YG��U��{k��L�Q��$'�a`�PF&Geϋ<��<¾���y%��<P��XC��5W��w-'���YqN�L�d_��r#
���;،��歿Ԋ=6F�����>�)�u�zQ`�%0W�X@���Rʛ��R�d�Q��Am�Y!�4�\��J���r�(0u���<p�����h4�f��|�JY%Z��&L}�i�m�(S!��JA�ET�i���=��{�>�������8��/��7�Q��^�
���W10e�{�|���ۛoC�^�A���G�|;^�ܣQ�㛍�s:[־7w�T"�f����N������9��$��JI�I�D����|�Kg��n~̀�0����Z����Y�̇߄}V�yh��k�� ������~݄��(�y�X�(�WD����6\��[�u��<z=�K�ʎi�Y�w�aO�i�B�$&�y���VAz��u:L�����A%R�}��E��hlZ�d�A��F�D�e��q�{]��39������	�2��|kDrӝa`�v��H����q|K���/,�񾟸�7R=4�$^#�	�8=Tqt����쵘,X�v���ڽ⨉���u��&��z�G=4h4��L�yP/RD�TCwPA�]��`��J�2%�n�d�_�ϗ��y@�C��R���,�-_���I9���d���|�ϐ�V���`EK�n(�G�֎	��P�z��&a�h6� jo�߾�yx۩�K'M�����
�_t9�t��t�����	�u������}���T�L�w���ϸ��ǰ8��MƔ��8��3��s���Eq�_1��0�9�Sd�1KP��]�<]�;Z�u�1%�J����,�\_�!���Y�P�\�r.��2-eL	��5��M�@魂Hcs�?;�R�$��|�D3���(Q�sMS��g*qO��I-b�,K\*.�M����
L�6��6,�ϼ+JTrh��M ���$������/X�ffWL"o�'f:ǘP5���J�T�� ��D
����<����x�_��;Rg+[��É��]-��[6��;���T���x�]��	�2������ݭ
�3�P�b�iN~��qﳞ�w���R,�7��#�eq��샀R�+Ղ��Sl���������h��'���p:�L�P��>�#� zJA��$�28S�_:��À@$�V͏���� rՒLc��R����ԟKq3}��pe���N����ci:Ӓ.��<��&�T�e��)�1i��1����kŬl��j�9^��\��#d¶��Ɔ�f�f�2��!�t����9aI�1tCzOT���RPΧuGbv߹�9�@��h{�zmq�5�ХP��%���R�v �3-�u[�N�����W��x���<+��X�ʠ;���\�{i���%��.h,�*�h���ڍ�����fLG�e���b��py�!7��s�t]O��t^}�uk�	�W)��=g�$��!B��3��;_���j嬮I·w���O��~���I˽t�C�x�v�����P�5B����R|䥱@"_֣�=O��L�X�a?�o�����O�ب�<�1���7)r�e�`ګ7О߃|�@��F��@a�"
�O(3��.?,�HF�q/=83��L��3eD���E9e�n�/g�)9��S,���Y�B�(�5�
c���)���[��p&q�ve�H!?g=�,Zj��6 >k���4G�#��Ɣ����K�CW^���"Bk�c�1�~�V�O���Hy9���ʈ%��+'qw�h-�v���2��V�ٗ3Ù���7V��Z ��Qd`����B&Q$��d�e�����B=Q���(�z�2L����A&���3�O�߀)����ݺq	���%��[E^xȁk��7��:�h	��i���o��ގ^���Z�y����w�	GmX�#L
�Z)�I�=C�9��ӕ7�U��\�	߽�j<���R��0rTDaw�=z����a5]�M�{�M����_�G��t�XܽcU�M'���������U������%�����ڕcr����G�z�8�'c��qI�[�,��p_9�:lz��\��N�+	;��j�sV����1�Hv�R+�X+��Sn2��Iv��^���%��}{4?0�[�$�Le�jlEm�]d�ELT"컲�U35����,�9lߺ�sduS�\�P��;���yG2b f������TtJg:a5G*oC,��{�)���x�K~0ǕK�Ǧ���@�@�1
������
L�؂�D��S�jR��ص�E#�bg3L�Tf��1�aN���؎)0\qM�jE������Մ�#8����uȦryv�4�u���?ԍR���Ŵ���g��՞$>wp�֤�Ӡ7�������"ǂIؽ|��?���p/�~�FG�\�>��ۦ��r��E��mo9�_B� lk?��~��][�ɍ��(pޕ���_�VW��ܒӕ+��Ɣ�T��ĀK�JW��h�:�,4��W��7=���q��4?�۲��7#Z�[5?Z�VY͏Ls
L�?d3�3T��	#�r�V�gH�42�f9����R�b� �
����4A�^�#b��T[s"��1���p�t��~�m�æ}-�����Wda��}�z}�K/��v-b��r�Z�k�Y-�>���ٳ��E���5�9�.ep+�*֮[��fQ�U����]�v���`a~l����d<��YYw���젛�	\s���?c��3x�kO��3���:�ah~t�ߝ��"&W���r)4p,+�Ri7Wۘ�bO]]�J�R� d,�j�i*W��L��9*��8!a��;�XY�51ErH
N^0K�lG�!���(����L��[I���$�t��$��f|$냋c�ݡXeb�Ӷ��l�=���]q��7��ˇhr.�L�7��U0�*��߈�! �_�V���,a�<�ϴ8/1 bli<�ƮWb�]�??�������]]=8�����A��Er��0�U�4)��O�]���l5��d���V=������~9׌�##��DD9�&#K���(`,�^�J��u+�q�!`��زc��>:�^f�|E�������^,\�gk�!�� S?����T�u^
ch.}�'�OǤ	�M%���ӀɊGZ�V_	ieq^���|q���kA��|�s�Y3��-���"��S|��JǞt,Y�i��[��"�ɟF���HɮE.l��k R���~&~�D��-y޺nc@g���j��\?[�8��Q����D�����g<	O=|=�OVQ#��K=��^O���h�E�b��ݸ���p�a��z�MI+�(k�y�B:�]^��U��,[6�v/��6nÃ��0(N���\$��oV���f�J<�h�0���<�|��M�#dWF�J`'&�7L�݊�����x��
� �BAS�Ű��ߜr ��M�9D2GԔPNP0�d!����ZX�Rz�ќ���羗g	Hv5�}A^7>��g���"j���R�g�"�B�, �c(�C����Ctl�<s$%�"�=��i��{�3�O8ǔ������������:`��֓���jQ��7nY���#�p�m,������'����:�;�D�T�\퇺ET=�����\8��[p��w`���H]oi��j/!��Ƴ��_��{c`���ݼ��͟a��,�ކ�� �z˫��3^N����^_~��6^���j�$� �}��q�߉�؇q�	���A��k�����خ�B��tS�s4��"TT��:9`�(�=�t��NIF�Ħd:f�	����&h�׷��Lh�AT�f�ܰ
=�M��T�����o�9�\��;��O;]yɜڐnY�>��eA9���.I҇��̷n��8��t��{�����zP|���s<��^y�$�M%�,"࣑Ř��Y5�SN~:p=ff��\)����l�9���M��Ʈf�{���WȊ2�!r��qM�@� b��
��d<%�V���72�Fz�'Px+kEz�	h(9�����D~�17�E`�ssUʡ3^xZl��4(W��{(�s�6�0U	qġ`���m��y��-5Y���
��a��-���`j�r��@<��+�e��M�ꘋ*@e�0�]FY��E��ⶺh�-	0�~r�j�'�pFr�èS픤|��6z�MaL�=�ڈ�F����/�y��I&P���H��J%2@w~������3�l+q��a(;�z/Ȍs���)%-��,NF�=�H�T-��e�����g��"��E�9�Q�Q���C��Ao���!�C|�3�0-�~�|�Y���QL�#�r�f������Ώp��J�[�T09=�b���2X���bAL�K�ɑo)`B�T��{�)��4�v�h7����z�r�����㞁��*Jt	����M;p�u7a���x�ч���~=֯��}����s�g}�[���0��@d�ҫ�I0�Q��'��dwhpԳ�����,��9���	�'�s/(:$�4%�4��P���f�%Mu�%F`ym�M�X�6`*��Xy����=���=e��ή�K�R�I�^���?��F~�Lf;�|��Q�'G��=Nc�3�-��ǸH�j�E�7Mz�8�=����mf����(�罏	�=&���DP�H���y�ܞ����1��sv��'������2H�S
�z���dVMd�� ſ�Qvnz� V��B�-k��� ?�g�CT���#?'���X�̜�g>�/Kg!B���{t�:CjĊ��$�%�U\�1�*t	k�{RTI_l�v0��ޗ���"q��$�Cق>+��tٳ���oۘ�U�I2�$�`y~L}_���.�O�*�Z41��*�^yz���I*��E�fg�_���̈��-R|���Lz���w��xZaGׂ2{���?��������=ڳ�����'�u)����:�����[�X��c6���^�"<��M�%�aMu��pR����ѽ[��q�wb�6�Lр�HTk���#���³�Y���ރ^l|��ׯ���F�8n�*x�hq'���W�	y�^���@w2����{̘yz.�~џ��Gc5i!��{�\���ǔ�4'�N}�gr,�@���T%2�}zU��_$����E|Ν.:���
��*cZ� S.
H�QV�
L6�F�U��$���Q,�ӭ���o�~���Q�6�/{p�AO݂�:��>����&���,=�OL{L��h�^t����-,�+�{�v� �JA]I7m[�����?oC��b�����8�YG�_�Ry�:��_��z��V�9�y�����B���8�G���GЋ
�}����VkA{�?f?|������͏�_�[v�E.�4��>N?���{_.�)Ѵf۞%t�]�]5#�y. ~|�/��|��^�ib �u�k�k.��عT�c�;�	.)��~Q&(�g��|�R�RA$=>���){eCaM)�˰�Y�d!��مWptxm���S�"�{ځ���^�1�|N� ����|�����e��G`Jb��W&@Y�E��{S�h%�ap*��@W�БCr��7T1��p����k�z��Ϫ8E�>�d�@����V��ñ��>2:�������#�?p��k����π2 �y8��~+���/"[��	0�:WW~b#1Op��No��[�0�����K��<^�#��l4�j6�i��W����ִ�fL��׬O�O�BJFe]�AO��jB�!����e�-�R�b�R��ȹLaؖ�ߺ{�l�ڤ��R	ũ	��'���SV��l�D�hh�!0]� 9�fr�c�(奌��j���z%��(�a���x>sy�&'PZ>&R�.�J������,S�� �=�`�'@^̏hP����y��ɐ��1�"����,0�XB��>aI�3y+��=��0���Rp��P̧�9Ǵ�E�?��}|���,��z����f��K~��n���+�צ��`���ظ�!<��cz}9���K�*cc(WjD����\�,}��R��Mxln)�TH��Nc��=�G-D�*�ff��l3��s�DX�����h�Q)q�3����;q��3�wY������<�1,��`dJ㈤�Sk�&�y����Q
-�����N���}5�(b�D���\H�%SkqɓM(���s��u�oO�$ws�E -39s�E���ӋqT��{$�-�T�l��{F�j�0l���;��5U��i`�d���1�x�u�8~�f��1\�z�@�&C��Y�t</�(�Fq	��='�Ð(&Q�$LWr���/%�/������1"�"��ڏ���9(������ ;)m96�S��6��%�#�#��<=�uc�"n�ל��׸���Z�$1�������1��vug�~�,L򪰽����*mO�9��g���POzÇ�B��Zt\2�����8��/� (55f�-w���$� ��8���*�,���e��)g��Xnً+۴���t���N��ʼ?�Y�ڒG,NH]�J46$&=^�r�T�Sq��א6��<�z�-%BY��%?�dp�j�^\��`O�'��.��3첨���Z���X�xޓqګ��'�GYz[���O�/Dq`s�ů�&D�k��Ww���+l|h�r�� �>�@|��ހ�V�H��/��&��o���P��r[pd���Gj.)����X&����	��g���~Ɣ��2.Ff��GE�<Y��    IDAT��g3(q�Q~_o!\j��f.�9{L�r�jY�Ki~$�-+rj�A�!'�f�:��;/I�E�\Fv��l�(�kS�����#�l�^���F[ j6�z��HE%����g���E��Q9���$ߨ+ui~� Sv�?���)ݢ] �����Ǘ_�m;w��}	LO��N|*�u�}`[_:�'��7w r��D1�pZ@����1x�	����c��)`�4�0�v�����غs�<��v�q�C;���i�$�t�d������}�8�s�Ê1E�쏸������z	�l�y��=(�{x�k��O~�dL�rb�{^�����^�[n��/6����ټ/�����j#.��v,���S#V!�^�V[X9��%������;.��9@�Q�t@�,V���4��/�S�#*6�r�p���Bg2��,GŴq�!������t�6���7���4Z�4�i��{�R���U������00��Tn,i��*�`yp���Ç�����>��Ƣ��hR�R
?<!R��{��@�_)������5�	[����ԧ���|�-׊�b:e,��,�����w���VTB���Yieo�jF+��P��KMJӒqB<�T1��\;em�{���?K�m�fKf���챨A�(gv2a�Ti3�4�}��<hM~"v�d�u�3����^e/e�ĳ�y(:`�ܓ?��0~������G�2	T��O�P�"[���~�����T�����{-aLs�X�J�iXB�Į��.�Ä��;D�6��&�6����(W@i��t\�i��s��;�9���m���{�6g�*�S��%05�iF� z�9��}�1����.t���u�g06�SY�����_�u�I�Оφ�f�p����wa�zL�"�9��߽�^�{Tǖ�69�F������h�^uie/p�T����9�Ƨ�99��tDH�����*K�M����w4wa6��Eb���.&��J�Z&/�q��4�q������I��q1W\��t!��>#W�G^�)r��TRR/��K mia�K��G��άKT�_�2qHu�T{Ʉ=M9�jL�yt������R��8&���&<��7N��sm��
�e���7Y�ƪh�!Ce�Z|����{�Xhl��.���M%�qQR�H4텂Sq��n�fybiYd����&l۔i���RGa��d�sJ�
ݓÿ�fN��]�3(�rǹ�#O$�@�S��uǷiCgJ�O�'���/���5�e��Z�2ɦ���Md1c�����wd�y��Ł�;2M��_7Er��$E$�nW�qja�bi��f������"������&��d]z�^���ǜ�g�_��?-d�����KD~�
Fޏ�*%u��5���B���v�>'��AgR@H?G��d��W��zp�g�׶��~�fNV�1%���e�ʆ�v*�yUO����%����6�3��ܝ��ilN5SԄ�"x6�f��N���I���>�8�8t����<���/�R�3i��b�� `�	\q�}�׳�]sK��Y���S�����NМP��==༟܍o��FD�e2�*69'���\���C#�R7$�?SN��c�N�4?��c5�R�7a�<U[�*���m�E���%�+aA�&O�����ʫj�a&ۼFXl礐 Dgq	Qۀ)�ѕ���V�fܨR^=n��0I���(r*A4@��Š�&�E���,���rE�R�e�1�K�^���e/lH_� ���7)�akJ������6p�7�K�Ɩ�۱��ex��߀���0�no��s��{'�Q	�3�E�j̣���)��(�p�~�𴣎�a��eS�P��#���`��ݸg�C�յ7a��%����"�P9&�Y��V��cWz�:���܆�y����a�� ӫ��!|����֦ �^{	���gu >���㰃���5�?����7��ٌ׼�%8��8�"~���s�/�������j��T&�|��H���cc�r���l�8��P���A��eʀ��t��5�d�g��U�}����~�~���Z!�X����Ȼp���A��o�]�����c�I�$�:�D���C�ԥ)Z������Ҝ��`$t�+����'R��It�LO����װ'S�Ϫ�K1~ ��fY�������@�)��~�X�r9
E��̵R�5 ��#|�'�æ:�"����j߅w��M�8����/@���Y�2_U�<@4y0��%3��v��f�)�qYܠP��Um)26��\k:�k��M����!���E�@f��kg���'ކ��	۾s	��9��������'���lR]��C/$�2�x� �A�����-�؃����|��+��P`��P���	���ˑ�t�,d����)� S	�
L�3��X83`�[�~%�w�[���Z�搣ɐ���sy��
c*�XI/��6�-�
֫�D �|�{�%B��blU��X�� tv��k3Z�0d�;˷�aU_���)+@O�عk	�m�4"�y��Cֵ�EJ(����5����������z��$�\Y��)eFO�d�k(ٔ���ײ=�v/<��X>U�-���_����/���Ru�s��1�|+f��f�0�zg3������~����;�bU�I+�
L^Su�$=>A{�=Y�G��+]�2���^�8PƖ�}��埖奀%�g9e�鐙��Ҹ�3�*iQ#�T�(�����◎��k���;��;�k��kΤ��s�:&K������F�Jgk�����VJ˅�i�
Z�1U�����+�1�1<�3�.x�C�rC�&q�2%�����>�@�kK�'f�� ԣQO,��Cb����&�U��|�cL8B_g�ة���5R�%��仛;h|�)Q�ݭ����!z�����Q�B�gɖ*�U��>g]�o��n{Q��o*��3هɽ��^�zcm��}���M����*��D9�iV݋|��]b^�iv%���=s��
��5��1��mNמ#����Ih,�"e��9Y���P�v�uu��xĈ=G�/�.����+OH�O,�=�e�2�{��%��}Ǒx"���M�o\b���c�GD1�^�n����E���̷�V%������S���.L��Xv�|>�PBnqDz �э�������4������O�HF�t2�c��>un۸ �)�~�����)s`)����p찵k�?6w�_��9>���P@q|L��xC+0��&�
�m������ouԸ�9	S��ժ�-�� ���[5˔v+��_�-PA�!��R4��#m��l��n�]�����$~�T(]���r�y�D
5��7�leTМ���TN8>o����a>�X�E*������.���b"����^r#.��Uز}�_7#���'�r^%X�_�֥�ᦻ�A�S�����/	m>
��Z��KT+%T8��� �ݛ��������V�����>��Jb�΄��@):����܆��'{(��ܻ0M��j\}�C����M�CH�m{��x�1�����c�ހ}�΢Jp����^��_�[d
E��y������(�����q�/o���nCֆ�k:CI��B�C"7VQojUJ�䲀�ؙE�TD�¾S����΄�2@�|�AY�T����$�|[�n�g�zu��8��Y�~5�ղ���7�ȈV��\��fz� r^��~k�Ӑ�2�8)�c���S��p������O���xi�O'/?���JW�%����W�}��3���r=����i?`�_2[�C�1O;
�l8���gZ��z��K��������Vюh|�k���x�%O�mYB����-�)�G�Ww3M�<Q�Q&������$�r���0U����D�@e�6�T�x�R��KS�񎎧���ÞN�±:�m�Ю�#5������z)������Ͽ����P�]���,��S����&ս��������N��v���D�TAuv���T;pX��b��([JW^��fG����&��\�)5?��,h���a��*Sc�H����݉��3�,��v߅1	�����v�b�g\�S������QSKj�o&U�>��̕T����L$��&Z4�j�&���/���1kc���V]s��%��N�r�r	�&�V���p�����^	a��A���<Ԩ"]��(u0��❧�
'�|*Za(��7	s&���r4��Z��>i��K����ha���A�,���H�,�5,�}���]����U��F6?T�v1�!��`4*�z�4������Vd�{���{��f��f6�[��1��Y�!���y����f�<i�<M��QSq�0��YC_���1`��t��$���z���0�0���V|�4QA��ad�(d!X<���%���ٰ����A������e�~&�؟� C���[|��� \�ɏ��(����{Z����p�-�	ؔ/)�J���;��0�l���Y,kӊ\
��?B�%?�X8SѸ�yy�RT�3/�Ԃy<T�M"��8��2N>/�	�d�}w]^*���*�8LW �g�f�+e�#}�i�S5m�קs��Z�{j��ď���H0l�  `0�x����.��s$��-i�*)�]�?1�_[��Mv��=6v��Z|9v����H�Q)(������z��S�k�4��E����^���\1�y���mq���{~N@3�6:��8t�q|��o�����8aJ5��{�ǌy:�,˥A����o}�l�`���z��Xs�£KlR�r���������`av�r�LN@�%����bLG}Ff;&�}��/w]ݬHy�2� ����5�c^�,��7� 0�l��NF����D���Z(�B�l�̫I���/�id�VK��, U��V�n�~�c׌�p��<��t2@����=D��:T���H��)���q��44�1h��E-Z�q&������,�όi8�d�,v�.�	����عk�w��S�r���Zw��s�n���l�
at�P��?{=�&��eQ�cU_��l��y��J2��nZA?�l�(��20[�qd2h�"cN@��:�[���E��/~�tL��t��s��_�o]��;�*�";u�X؊j��CZ��u0�xʫp��u��������w�ߍ��ir�~x�	���K�������ތn��A?�B�"=Z�J�ˡD#V"���ߝ�J�pg�&��yNl.tk�A�j����x�zr.�c$.^�-�����l�@1���T�U&�})���:z*����G���b	8��L��I���,�f|���=��T�K�9�0ؼ�������L��ב�?�������x�#�EP��6�(�AH��~�2�k� ���ͮĲ��ȕ���ض��m�u+��&�X����,�;��Y��!��T����d�S��T�Tӟ��H<�KvK����3���g��d�6�s����`" �����r*���u��v87G�X��BФ�`o:�xכ�%�ټ�� ��y������}��Z���8�qd�W�� �GBp:P�������ba�/WQ�]���8�B��Ԋ� +�칦��=��6ڲ/X�퐥c�qzȐ�BV�84�����b_{Hyŕ7Dwς�1��g[*C���{}�����$7l������6[�� K�Kʤ.< c�՘GM�#�(g���d�o~�,�?�=�NrؖJI�65�Mt͛<7dю�������x��1D�x���R;��/��]��	�bz��q��6�j�qn�'����s-W��T-n������_��h�+�E?G��u�ʞ9�j�bN��
�k�fYb��jb���T����6V�wʁ��
j?h�lY?�V�G�j�ΩB&U	�~B���������
|c��s闶��/]
!��9�'�]��d�gM��F�.g������D�Gf��0�U������Oj��q����Y'� ����Ybg.�{��wrH��aV�����dN�J��b��ܨ_\�� �t?�m�,�Y�1 �:S2Jc�e}�����](�`0�69������<G9�� A��N+�����@��]�67U��<k{�/Oq���jc���V69�9Vu��q�*��D|�[0H�t�D_f 1�DS� ����o�: 6i�������G;���#���u�2�/�Q�Z:�1�j		�8@0�Ϝ�������{�_�&�%kQ���sg{=�J�#���E�yI\P0�l�}�<,1Ƣ�P|<�J�^����7>M|d���v�lO�z����~<�m7�]�5��J�,�M��)Oڀ}WO�d}�<��8դ�"���U�� ����N|�{�ね-�q�U�e�Ys�9�j�Wc^;c2D��.[_Q"ogJ�}I`:F���6�OU�#�X|.�4Z�.�S�t ��REnl�r	�o���}�r���CyOZm��h�I����r�GZ�Ǆ*��CC��k�峕�����y�SDc%���c�(�)�U8�����a���j� R�O��ذ� ���3ë�>��h�E���E?�	����ع{N����/9�H�b�>�����}9n��N`P���\q#�w������b�<�>g�ЩTQ>��(C�LW`�$�:h������Tܟr�<�&"uԛ�1�����?��ɷ`�b#���!|��_`�i�~-&�
�.ڋ��jy'<�H�������{m����=��j�]u���m�?�n��fd
�S6����\.)i�I"G�Δ,���W �A�E��;�ߧ�g���L3I��9%�E9e��3iF��L����h#�o"����}��zŔ$��F�w����W�U��uT��'����V͏xy>����3�2���P0O
�kˀ����*�� 6"d���l��U����$̑t��y��P�*0�Ԁ��;��>���8�cS2�����+��Ǡ�
�2��)�bo(�j�r����ڨ�o��E �J���a�Z��&;u�
*��T�(���V�"�D� ~�i���\FHa�ó��2�1��k�	��a(�d	L|��A�|�����~:*�g���,ξ���w/Gi�~(L�ByvP��V�~r	[`L?U�N�;v�Uo�X��23��8G���7��&0e����ba����m�0%c*�����q�g�0(��v�|}�s���f�F;`�k�P�D����r��c�:k̊� ����!�g.���@A�}�T��R !�0#@�/�������C�E�%����z+�=b\�d4F8+�2�H��hy�<u~b+�	����
�d�t0�MY��}�Z�3��>��7/�_�T1Y�1�5�%��0�m�̣
5��6�Q}>����Obv�z����l��@��/$�4���M�Ś
ERvgLS	�+��ђ ���Y�-�%��8�s=4V �np,	��j�]R�U<�^��(�f$�|+��V,�=��`��&��00b��G�◯�1��;0U�}Ξ��i�'Ö��ܝ�9��&a�'¸\� ��Qm��00MV���b��+c���^�}b=�L��tvQ��Ηv�7,Ō�P��V)-#����?�� 9ߤ�S!��9���է?���Z�A(��ZG�y��F���]�hc����z�8;�S hN��!���֒������A����A�/*+:흥a��p�>�%:��XJA���,��ٟ��Zp�W��x�0W�����'aA�+��?]�oI��͍�G�H����zH}�_1�.M��|+b�sq��|^2V����P�ܵ� Fh�(������'E�����{ŘیqN�c���@��)�|� =X�^�A��.�x������$'��b�3���\��y?���ߌ=m���¼UϜ�j	��_����<��O������ⰲ�ǜ��1T��P�^������ԀB}*5s�>&�
S�rmd�@NC=�/0�s�u/Ym�Jr|�rY̗$7��+ᦳ��H�H�4;��/��T�B}�5 *ɥ��>!ޞb1�䄵OeHV1/쇒��VX.#���y-3���2�m��G�}��!e� �    IDAT�CR��p�����)�I��T�L������xש���4�G�n&�G����5�����{N����k�x=d�q��?���gd%̒Q�s,�|���^�����t��NL�d�׬��%�T��q�q2�A���ӡ��A�D���p7^�����<L[}��k��߽
�l��n;�%�
�veG�'{��]]9]R'L&Kl�6�-���� ���[���n���F/�� �"ݭD����J�,�:�ٳ�����J��dA2�qN#,� �D�&,V%C���hb��A��8��D����rh!�1Y	�y�>�`LM��l�p���p�u7�{7�h���Y�KKS.}2��
�`i2��J��}�ށǕ4�2�td,�UK�����Yr�$�+��w��&�g?PS�Tr8��� +͏}��uE&�~�}p��c���cl|J� S�������l�-w>�nq�┍Pw4}�������:dL݅����ߗ U"\4�bFđ!RtԽ#1�@����'YJ{�~�#�v�\�,���d��N��u��W���0���Tp��ʅ�������ǐ���w� @���7�`�-��g�/߻�^|-
S�"?��ٕ�T�dɽ�,7�{�}�"�N�;w����B���,
cc��/�AS6=���U����F��������ϩ��$�%�R�L�1�r`�e��7��l�c����2�,��	I�2*	VʴʽS�:z�[Bbn�#D l��$��_�kW��I��O�7Y�B���8���W=����E�J�$gIy��YbY���%��	7Z!����_<�n���qf�E?�nq?�t�M���
}���c�7?3��s��Qw����� T�]��(2IX����-8�?nD#�bz�:��S}����(������H]�@j���R�p��f�c��b��_Q*kRLK(�-O$�r�J��=��Y���%o����2�K��	{�W�1��9;e�,���تE'-j�Z��P�'��<��_.31��]������Si��P�q�Έx�U�5e��%*is`*�{!Ye�,����G���ۋe�iH�?SM��T�9Z�4��V)&����]o�<�G8�H={?`�s����L����
����2�����z2vT����	��Z�^J�k�ہ���$����5���CƼHd�۪1��N�A��"���Lf�[1�thʺ0s�����['%fQ�mN䲾Gb�i`_��*�z{��ڝ�=u���9��d����9�lR�JQ�$�I��I)�-V�����{��G�s����}���{�Xr��bb���<n(�K���ev��:�^�3�yɍ��ܸ�jJi6\ª�>��S�cW`�k�3@C&b܌o}�l�k���a�"�&�,}�U��8���������k����bQ��6O����/�{)�p�f��32d�U�CO��n*�S��%�qq΋��*`�}��q]���SZ�H�)_�9��B�r���R�rz s� ����X����f(�%[*}�t}���2PaI��~��ɲN[e�\��"
�
b�D	����x��`�l�YoFLZ�����w�c�<�B2sO1�T`��z�Ex��3���N��+�7`:����m�����~�ť%��,�z���E�{2
����6��s~�w� ә�U��ʀ�8BBu��^5�aՅ��'0��usB��I��D�J@�Ü��¡5a��L�/?�I��Y��:%����<�/�J<���	?@���S�o=�$<�i�1UQ�.n
U8����K����XI�gu�8��נ��*b�L�:>�L�n�9��rəK!m�Ct� ���tՙS.�\� �j��.��ڌ@�/����=�b���O���J!@�v���wc�PvƲM��_݌�|�-����	�<��hЗ�c���<��0P�L;�R�����ox)T��U�aG����ͯCH�Xu7
.�2W�t@�~OV�"��ic��+�|��Vt	 ��׊����?���?��Цb�XҾ�WV���-X�I��y/��&I�53���(��ޣ>�v���9u��ň�;2��s�T�ug ����D,�����z�j�B���t��������Ϲ�A{�\g��5x��"�����S߸?��P�XT���b52���ګ.����Hb�'��6v�`�/�0N)��"��)��Yx�dB�@�K�@fr����W� S2���e����\?�HCzL���x)L�Xc��2)(XU\��7Xa*XHH8���������w����؜�c`*��3�Y'CF�;�⠁���`֯[��ZI�+t��z���7]�d�a�5L|9:�����a���6㷷nD��ȗ����^b��}*�nV�iXP��x���x�I�`�L�J�2= ��~I���[���E)`�IZ�H��V��W���:��b|�
�ÓRS�e�����h���N\ҫ�(�T�`�Qy�n	w���q ��l�v�l�G�s1c̛'C	(I�ߍ�i���Q[c�t(4���T�KQ����J��[q/Տ'��ML�K1ff2b��\�U��r6^�� �`\��e�j���Ԟ���K��]s�4>><������(ee���?��cD�≼�7Q@�n����T�3�㞀&}u�����s���L���Jj�# ����\��L09N�I��_�����5ųFs,ƀx��{������@��m�̜>��q6U�sß���~:�ͭP�T#��xE�x]�\su��58��*�rK�"S�o�酙�wK��f�WS�{� -/��|�f�zې=�W�Z[-V(ӟ׼7qg�¤n�$��|&ub�E���g��%�d]�i`:ZH�tY>2�k��x�w�H�s��V��9�m�n�H��k5��v����4������Frv�e~�m.¿~�Ǹ�w�J(��l��R���O����`��|���K�?LJyl�5#��D� ش9�׾w	n�s+��2�\���Ų�I���(=��-�ݮE	/�H;���ϒ����Y�rF�4=�JED2P�wRG�9��\޶ı,�R�fK'.���I�LV*2�T7-�����K�r �x��5�ݖߔ��'ǰ����ȄyO/��N������w�-�� ��d��@?)��t;��Q�~�h'0=���R^�@w=�ŷ.�W^�;,ԗp�����o�I��bv��1�g�{9n�ݽ�c:;�Jw������:I�s:���]�M����~2P��?k�A��H�յ�0��s�� �W��|�נf;�=����~|��+�}OO���:�'�8�9G��g����tƏ�K!�e�<۾S���f�Oav��5$�.^��k	���a�GM�$����L����+�(�A�+~Ոr���j��µ�XV���C��R�R��c����p��L@YcF���"Jٶ ��VW�=�'�q1�.p����/�l9�xB٧I;-s��{�K��Yʔ1A�P��JB;�c�:q�;������14�����jhr%q�v��H��3	���&��<)1?�!��n�,>���`��"qu�li� � ���p�͛���e�)���irs�{���X��o�K�E?���H��((���!]�&L�v��N���t��!��?eK��X��z��0���˞�D�ѐ@YM���zQO��+�sE	��<�����x�[_��N=F��x��}��~-.��(O�j�P�Y�L��T��	���� �laq�,�/ȁ3�j���F�K$5	�\"7h$�bSaK�
L���P�<9����א�3cLy�%9�������/���d}}:�G���*.�b���L֞�&����zL��u�T4��ⳏ��%.��Wf���f�<2(��#��;,�Q���@-d�*Al>��ř1O����^�a�I����YV�'�B�BE�,QLh�B�ߨ�"{���a�A��b��B�����B>B^�,E�_Z+�.#Ty-�[r��dD�~a��14���qr()f�$ӌ����pe�2>&�󁇞9gz�تѲ�����6mX�̵�����d�ɬhs�He����$xGd�B Ơ�c���ϥ��Q�T�Y�q�5��%aLS<��{�+��Dj�*::+����
���V�lDK��pJ%�
�T��s%Nʼ��{�4�)89$�XSEj��:8��M����K��u\Q������.�H%ǡCM�7�Z����4U<��U��3�$��_ԡT ��w�E�~���KO�$���V�U��R����#`Dg`{?���&|Rv1�M�i�^t���s+hXQZ�(e�g�+@��t���6�d����	�ij�0�j\v���;�3��[ܯ�z�����u�($[0C�C�?�>:5;�<"�.���<p`��<����@����K��Ѝξ�$�$�K�m�-ɺ�U���Y�|;�����z�뾓7Տ�U'4|��^�����t��W1[n�3|^z�:T��o������E|���M�GeL̬Eu|Z�e>�A�>�������4؍�;��xӫ����
���"���F�C��貛q�o�D33�6x����BZ�L��3�՘L���`'��b�J<���AL�e��&3b�G`Z��E3������B��T���8��@�#��޹<�r��qd��!*��0�B��O6��\8@��-U��A+��4P�8�r4
M�����>��&<�q�����f(@UU���q�� �
Lk}gLO�3��E�;��b��H��������cai	�
>�x�����.�P7nmiv�� �$)�^~:�yc�J׼�FzKe�����O���k����kY��:�+Mt�$�Tz;��_�)�#{�.��^|�;�Ķ�]z��=�^V��_�|�����qp��o��.���a�_	��ĸ��c�~$^��W`��G�NĻ�3?���pQa����d|e�4gQȪG۔����K���~���%Aʣ\.��0�:OxyqDF�b�YF��M���\ǲ���O��U1H�}`a��_�K.�Qh���I�*e��Yr��Nm�m~�k��W�����|./K1���uLk�1p�^?��0U}���Vy��Np��I��ø��Ɛ����0�s��+�M��:p?-b9Ơ�ľ 7ݾ��f#v�
聳�؟�ca���� p(�:l��3�[>#Q��K�b�D�<'�G�c�k�>�NҩY��'������e����}�?vB�mc�ߛ��|�}k]d����ٮ�W�w	",�G�
�?g��嘞L��?�}-~|��06�/
�3(-�g0EY:TRz��`l�1�]���mC}n�J3kס4>���5s���OeEH�Y2�\C�]VN��ÀX�(c:=�����hQ����yo�����\/BonA�q�zĀ�z�$Upd̚0�j�'~�&ISeL��Ғ\�,�ss��\%^�(�fYV4�>�e�Yi�̼� h7Э/"���ڳ!��$��i�Ϊ*��Ȅ9�[�l肜/TI�T�@�D�ee��f E+�����4�+��Z�-��w���A��(h��.�dxUq�@Q���6)���&�\�ೌbu�R��W �+#W*�U7�b�F�(re���P��_(K�v���T��ٔks����s�qA,
�jJ��R�2�sD"����8qNI�bW]W���5N�FVQ�U�uX�`���33NY�]�;�ȧ���z�x���d��dؾ����X-��鮹KK��2hkUPE�<
Bo[1���%?kb3 �W���(�pCs���i�0�9$3�@�	���+��W���m5��WJ�0r;4�����q���	i�>����2R�����Ɩ�Y$�㥆;,�q�� ��J93d-�h#�ͤ�&)�b�s�TxcM�/_�}<��G�"�>�	�?��0���>w�z��x�4}?���.F;��Y{6ӿ�E�X�T<��MN�+�EeFmu�,i��s�XO�7Hȱ�GH��{��/��u�ص&�ALϋFS���%2�0e�h�ܟa�H/�hX1`��W]�bɳ�+g��m@D�['zȡ�s���B������?s����=@5�ݵ����Ȯ>���ȏ-C�6.�0�6����v<v?J�]��|=N��0QL�)W��Р<�h��.�
7����r,0.UE�&����ʔ:+/����l�90��R�+?<$��1���R�H/hDC�qS5?�:L�O����V �)0�I$S��t�S��������%�Y�󂰺��u�j��0OjD��l�b�)s�>��l�� �L)�ߏ9�����[�|Ʒ�н��׉l�0�?��qR��@Q�(0�����L�{*�/�9#��x;g����p�|�R\}��1=�������'��L-dq��:���W��[�G�_Ċ�1���d�d<�K�d�~�8����:�R7��@�5���C�Ԯ3�0h �x�IG�g�F���\z����w��ιP�i}q7V�,������0nX���k߼\t	�}�Ӡ0em������$�:b�,�mM��ߺ?��^��e(���KS�
���� )Pb(�TF��1�0��N<�D*�&}��R�J������LK��ՈN��~;D��F?�#7h!�Q+����;3L�s9ܿq����wσ(��>b�n��n�����E͂���T5�@>c#_�����z�t&��uI���0:6��W��у)�G�4x:�Ҏ�f~��-}6?B�Y�.�z�{p�3�.sj�2Ș<w�L�����F#��	_$	|�8�}j�i��N�¦��K`�b	����f�2���z\�Zmy�l1K��LG{�ٷ̤�ja`;�8=3����ӱNa�LC���A�G��E}�#����f��r�A�w�U����.�ٵشc�镨άBy͏J��:1	�J+߀��A%n�f�۶�1?�J���5���:CWo����h��i�je(�f�^G�\��ʲ)��M��N��E��|a@��Z~$=��1kˈ+r��l�b,��"헐_��f�s/ �bL��$	s��;a�m�Y�2�M� S�K�xỶ_�ᖽ"��n�v3~�|��>o�	*{eXH����g�&��g2~��U
f���W��l~�|?��Q�A�C{iA�؏^+�;
%&@�`�xx����z�9�-�/#[� O��,��I/�W_��r��$O����R�9c�,��� =lb&Γ�%�^{�� , �]��Au�$QtxA̒Ty�NSǌ��p���5��Pf���H%O0E]dɱ��8Ί|����R��}g�7'c��x�m�՞ϡ(�#z�ƣ�fC�`&�d�t]ؾp`j,����z~�2�n�mE�5��*�.%�5�TKh1�m��f�S5~K+�0v�N.~V��d�h	�?�ר�\r�e]�V7�Ad(�q�A��Q���`t��cW�8NE�B���E�%ʔ%R����y}�����g&3\�a.���b��Y��~���IQg�R�(��?a�GW��v���kˏ�yh�&%O������O��>����-�I�g�u���>��Z�F�{l|�F���|�ݗV�����Z⴮;���	05�4N0}����L����4��q%�5{Iր"51Ռ�<U�����5�iב����?~��x��֢�m��N���|���a�c�1�\e�J	%�:�)"�����ο���������0^�SB'dk����wq��
�����d&1(N��m�J�T�C5 �\MVE�j7-y��?�qу�(q*1��{���Y��1u`�⧨Jx�{_;�6I4E�q$g��u���֞l�r�,H̷$Y�w	2sF���B�1���/���#��m5��ё�$8�Aͫ�TN���-�MK��e�!���L�9��!-��!�U/�1����K8���;O���2�}c���e���7����~�ko���Er�*|�����cB&��<���~�����";(a��5�|�����P���%d�R����#�r	f��pY�sl�y    IDAT%J-օ/	[�S��G��ZT-^����?�K߻{tC,-�ª55��m��;_�4�|y�����\�K�"IFt�-d�v�r|�_>�c�9\t껺�y?�#�w�o��N�<1.7]���t�K���`>+�l�B^@8��V�% C��"�`��I�Id�L�JI�)�@g���tu��e�Md���=L��g�2�[��b�>�6?��N&¼9��7M%��n�*?��1Cv.����T��2@qy��*qS��H���8ũ��!�	Y������'���T,�h��55:�u���ƆC�_�l8�P,�����D3�㑝\y��Ӧ9�U��8ȢT*k2.RC�ԋ3�2�����ws��3�[���C� -ѳ��j9ב&l���`�Oa �^�=
�l��� /��7��8�tb���I��c��'��[h7�h�;زu7�{#��4(#+p�����e��n��L�����Gqz�j}���� �Le�aq�4��0>>��իP����'�7gP%�"S��IRŤ�߿�l	0%8(�P]��e�b�Dy����˦	Ѕ�uCt��i4Q2���q1X-aK�(8�f���K����9�)��ͪ2�̼
���::�E:�-���^�J�2�2��Y1�C����"Ŧ<�(R���(o�I̚���H}�l��oRFa�ܵ�L�d�	å2���#@�9�<��D
<��D���Ѧ}�S2���)��'�2P�N
6r,�)s8਌#gy�yq�Ň��̓��K�w,R�,�����ʵ3� E5䞤�g���P�;q�d����^���r���S�4^~J�~s`y����˯��=di��ۆc�;p��TԵԚC�X`ߛ�5��6�Tk��Ĉ�׋9e�ч��~�b�h}��O��AS��N�+����N�״��1Fp�(ʢ�1�#�6�QI�ͤH)w��!e��g�>+9�-%���L�|5�����"3��ԘCP�G&h#���K��8���N�R�TJD��k�?���`3[�Q�f�8���d�
6�Y:Š;k���^�Ц�%��ۛ	}�g���`&ՙǓ�:��ئr��9�yl��V�ӣy�j3\7�����NS#؏�[xo���J[t���XZ��/�M�t��zH�hf{��C��3�v��/kq����[��9ޑ���P�ʹ�l���Q"��P��D�SG!ZĚZ�����G�AE �ɘ�~�<��W➇h���V�P�Q��Q���\����m�m8�-��{�x"�X���R�� �u����	���oP'�)Oc�1�c51���B��^N�5��R��< +���T�O�3��2O "�
ͅ�j�H���ǹb�,р�j�8%de�)�)M��v[�G��Z�\�-P}��bZı:�E�ꍕ8�g���o�A�2^����zy�+�����RV��~.��T��Y�[�.S#^:[<�O"�'����Yˁm%)�
� c�� ӏ��d����x 0�큦 ��~{;��:ݰ9�-x��`�A~d���/p����r��.g�$�L���B��l ��1��j��Ya�İC�_6Z�Y�Kbd�Gq�c%���:��x�IG�8��s\��W�	_��Z�䀹wi7ffK8���;O>�,$�����_��]~��؉^��01Y�1G�w��M2����[Z��܊\rZQՉ	Y�I��H��*�VA���i�T����fH�^=i���� �d�s��d��(R��F��{h.�#�,"3hJ�)M����@���jEX�
%t\|{��d����c�=�5-�����z�T��   Q� �bC�F�Q���(�&Fo�M�In��XQ,�BU�"���P��f��ӿ������>ߙI���0s����{����^{��6{��Hg��ǎ���ɓ!�rd�XŋH���^������H���!�W��L� 7�� |�`�WI��12'@���h5�Q_���RQU&'Q����0�E7UA}4���%sHes�K��A.�g�`F&u��e(�ʳP� �#����!W@�J}iD��t�e�\�=5�S%yO� ʪ�7�V#-��kZ[\c�a��g��~�+p̡:#ӕ���^?�c��q?��~/�}�Q<1W�bN�ny�<��2�*&�oDnz5�SS"�d�^�6SvO��D(������h/.aj��t�TE�YUeg��nOb�0Y��.,f�h�1m�Ѧs+���(��Đ�t4B��9��,J5	>� Gƴ=���2C�fb��B�;���%��3��u�	wM��(p'����"N�x��c4�E>3��wmO�m��I�P�Q�QP@�^,��e���ﲪ��EYa��2��X�u�CE
E���K���f'��v�y��F�x/E�7�b�%��~1ñx ����/4f�L�"��㽲����^���dT��1��j��n����rrdn#V�A�-�"_S+�L�q����og�zξm��1��Dһ"эeI8L.�-!���� r�Qv����"bg���!Ʉ�����2Q�l�(<AUJHy%�G⾮?�-R��١�\��E�.�0�(/b�hg��{cg�\�J���&�Y�2������cl��F��,��8OOV���369�}/�E'���5�,��]�>2�C�h�W�Ũ�O�XŉGn�������Q.�U�?Jaa��Gv��-w?�m��.�� _E/���?���5>c5�T�����>�2�^���?��!_Xtbɟ���B�`Ib������
_T0�?0�oH���5�k��E�[f��	���q�5Ի艏���=V\�b����W��3�������� ��g�r xa'��R�pMa�����d�1�0�~��wBD&���g���9vL���eF� L���\Sf�F7�n����+����L�*�*%1�a��ܾ}���0R�=x�[^����R�.)�s֍ʜ;�-㓟;�<��0���҅�E�4� ��ʚ�3(��Ҧ�%^�W$7�V��s�ƩB�S���4�S��c�՞G+$kO�"iɊ�4,�1	c�򲰦���kZ`J$�&g��65� I9�s-�e)���x�\r�.\�R\��l>g��b�4��]�l73�W-��l�"��]�@��i�Hp�υ�1�<�b~���7���~����X��&����翾E��S�ބO|�<��-��ZH�GL/�7އL��u�6�H��Y"ѓĲ��~pm��y*�wN��8׏}L| �����`�y��r���T9)W�C&�{�~��7�l�� ���る��1j��Q�wq�����z6Ϙ#�.�@�ݓ%��"�ݙB1�A��A�R w?����-���
ʓS:���jUEgjҐ�b�\���̝�X�n���AO-�g@���dN��Y���^��A��~����:� LU�������hs@o�-E .z��X¡�m��g�U�<�4�_\Us����ȝ����8�%�FB�����\�Iw�~�����c��21I�����K�^�&34��j�eJ�L�,��^�n��vf5�@vr#P`q"�l� ��������^'�u�`��yV�f@(xZ�=�!�+�X��u#sU�kl������D������������Ӗ,����^�:5���G�x16O�����!�n�)���ھ�܁[�z [�چ�F�|	�B�U����0ʗ1�˝�g����;�0E�����.-�Z*b��5�*�)���������$Y�@9
�3� �� S�nv��kQY�
���Yq���T[�c�����a�ZsH�����J�1v�d�#�*�>G[�'�.�C�jV��W����q�4]�R)j����5��B�SG��A�}�4z]�k�gVP�Z%}��}�7!�
]�8'��)�7>3_3Fپ��I5��y�g%ɶQ.U&�-���XhQ$ae���%��-�о���J%#N�wɚ $�uiɰ$�ξi�1�Ke��,���]������^�`�8�v��/([ʽe�i�H5O佚�]���f�ê��?�����1.�cA4*jE��HUM���ntӢdX��D��s�v&�����%�3�<��Ɏ� ��}cC5)�4ݙl�v�Y���rQ`:ξ��>���u�i��f9�LG�K��I��XO����G�P��צ�$���a��W���c�z��2
L��T����<�XzJu�$�{������u6NE�	����!���윅�������{y�Tyz�8��ߵ$�*��lC��hް��q�	�}z��=J@�ʢr�X�[䎬{Qs��ț��3���<�bs�Ӊ�UXWޚ�W(��Ic�V�S�=TB��c�F��/1L�Ox��r�E( ���l��	�ƍ�I}d,iĈ�[���S�O��T�����?�h�i.���h�f��v�R�l���sy^p�f���4h�z�͏���R<����F+V�L���0�����d��޷�>��XEۄ�O�;���|�]�'jUt0�!���򕒰�����F5]e���W��)�4r�]_���W��E�'�T�C�t]�[�,�E��.1�{�-[B�ؚ����iX��j�V֔.�l���N!G�J�JQ�#��#����uN�	sؕ��K�9��t0lҋG��r-$4h��6D���\X�i��Ѱ�d���%8����]�U�X�g6Ub��)��6�s�������k�ߊ��E����Gߍg��Y �;��\p��t�6"=��ʔ�ŵb����&J�����4'�����t^���0N���R-@��5(�T@�-���/a�ڍW������%KfȘ~���p�%[1WO��naan��9<������yN:z� Y����C;B�(Ѽ�>�����o� �R�I��Ud�yay\�)�Ot�*�d5(ͥ��%A_�k�H�&�z	2(㋥
�sy5RbE�T(HE���r���m<���p�3�œ6�A)��>��݇;�W_�+<�� ���җQ	6��+@�3`Q�a\-�ƣg��b���=Z��5Ti���k����������p^�>�p���yp6��ߗ�{y��9x#N8�8̬�6Y*G���a���m��\��~f
X�kHe�\z?��mHC����f��=e�̰�A�:ٝ�ڤ� �T��3���[��������� =堐��L
i��2��0PrL���ٽ";�)���J�%+��t��3�kp)�)��v�oSk���n�sv��\g�]-`8��t�T��7Ș��(���u�lci�^��NU�X�f5J���w�Z���2{�&�4�=/a��V��&��T׭Fq�$�ٌ�E����R���j0N#�!0�)oєH]���jEG=Ľpd��H6������n�,|�� ���<���#�ݷ�;�z��C���_�8�ux鋞���?J@Ƀ?�{܅�؍��t��3T\��#0�i�J����#�2"I�y���E��*alՁ�R���=I�]�����SY�ԩ�Gcd�J2��g��jZRW\�s�,�(��5��zIӬ�T�?��j��\L�������1�L�ҵ��婉��ΙԾUIR��mx�&�*\C���d�	�G?��˱օDr `�͟!n��,�PK�$z��H`�3�HC�q8Q�x��WU�E��ou�+�7S��C�}�]��ۊ&��YF��j�%�ˌ�΢�+�w�u�_��gV4^ݰ�I'����pN$�`�c�#�u��"I3�kN����m~�y��.ң.���������o{96�Y�Y��	i
�#1��ȍEಟߍ�\v_���A*W1�4)��Ta/�øY���;����4�K*�d�plX,'����4>���{�C��Q/��cU$d0�q�����?��Ҥ "�)=�I�����	 �4�IƸ���Kȃ�A!�^JL=ǋ�/�|+�`�qPC�1���&2��+��~̸0�_-hgcy���������ez��l��Q��M�ժ�ӫ#՝�!=��G���'(c�~�i4G���?������Î.ڃ2r�)�%*%)���K�i�܇�\�~�K��w�k&��8k6�]{�.|���G� mL"W�F�:�l�(>#2N2�D��GSA��9�D�P<�V,=c<芑�q�;�\���e	����d~'*T}ĕ� L�0�<f�fH&1��0�T�#��~����r/r�=E������9Q8fK���,pk��O��l�A������dD� s
��� +E�������8(��.�z�`>�'P�u���Kp���Ge��?9i3>������?ʘ�S�/�R\u�MX�/�)Gn�_0�$;��n�w/.��OqÍ�R�͛E:�s^�n�z-�����p���bY�#�)Ô�ŋ*[B�:-&2)�/W��Ez�Dn��3ZF�25j��O���y�)��'�Ek�!��Υ��{Wށ�v�F�ߎncS�>��mg�/{�8d-*��?9���n�L�o��Q���?���v�	�����^�P��8�m(�Kc]�*2M2h4UR�]Ta<��Z��ma�t�c\�#�`�� �ʇ�A�� O�\��^�<�Y-�)��K�Z߼�����Ő:s�Ӭ����g�&U3}��a8�`@a'�[���7� �̆j�f ��I`v�'"	�a�cG��_<��X��g%ѻ)�%�fZ�>��4�✷�/x��(��ғ�I/�K�ƻf�lŞe�&�A�~1�7Ʉ�2�� Li�#̃'�z�	�X=�U����V*b��瀲��t���.����%���Ҕ��F�Ь-��{]i���8�?�p�ak��?���Y���+��p�)��}-��˸���q����pv1�{(���u��}�q��1S�b���҇���j�D���%9s�e�|.�^mmh4�L[<]*�����z�:L���@���_*V�@�3@��i�)fL���2�_�
4��S����c*�Y�Z�5�~K�N���Ҡl�t���[���gdDUw�t�<>��/c玽8�Ik��~�r��}��>�{���G������� ��D6[�ă�jʒ������TYw�sy��A��Rh�ϊ�����*4�)޵��5.�!��Z�6��J�T����=�����ޫ��y�geɼ����	�%�&��� ��R�q9���d=?��Eܗ�qR��16�Gy��ST{ed�/n������x�����h&Hq���%�)�����L$���֝GVwE��sP�x:�k+����ö&�#�U�kY�#EgL"��%��
��7Z�;d�B���-^ax'=~l�rJW�$�o�J|ݖTQ�!�(�)�5� z��'���f���
}���TF�h+�;�򞆙����(�� �dGM��u<��u��;_��*{��;�lO��vX�2ҫGp��+nŅ?���*���r�pl�,�f�9hL��;��B�y#w�P��QC7]�.3�-Κ��;�e�Ozv�y΁��v�d[׀� ӡ@9a���t�&����+��>���@N?�- �ag� z-lyj"Or��FyTxsSwY\ճY�#�s��o��?L}�q�{�?�ϋ`~c�����c��|2R�0:B�R�^�� ��}�8㤍Ƙ��O�5L�ҟ݌��÷�k/�n���yW�!_*�YР�~����d��
<�5X;-�^V��������n�o��4���	�FaE� �b�˛�n��P��������B�V���	|��E-�`�{�y�ժ�yQ��(
bi�~�fD�4�Y�F�z�v[T���f<�R�K�V�/g�����|2F���<�d�4R�>�g�dX��{��m2��^=g=��mk��C�(E����UI�-ճR��x�Ӷ�s_���v͕���]\���pկn����;�|�w���o�[YG��;�/}�
��w�"�.����Ш/C�n�tk��8���p�1G��M�139���M�w���<􇝸��]�_ �	Tg։T�ULV�eq��-    IDAT�6����F�%�{�ڗ?���[��y>@�|��[qѥ���+ɦسk;�S�e�?��r�Sp�	�H�c��!��I�1ٌ}sK��q����,���®�41�t���s��	:�W�iGr���E�U�RI�������ۥ�hS@�0jb.�C3�ɟj���E��V�;��w�u:�9� ��V
0m���]�K.�Z�Sq$�&��`3J@����C��cK�4a�*Z"�1 �"	�Z�57:�T7fI�k�+�^ѕq��������
I�I��󔜋S-��3��'�
'�V��Ѕ	E*��xh� ]y+��@oDÉ���H!��dK��N���l�-U�T ���)lu��s=t�ֳ�9�E�%)��ŠE��v8t���=�����o�%HMK��;}4k��/=�Ճ�zx��i�|�a8��C�������%�d��0��P��*0� �x��_>�K��y�����OV�d�)�%0�߱��k׮���D�{�^_F�=�&)�祄7��SuQbG��B��Bˤ��W�03)���#�'8#k��:���;=�f�i6�ǔ��2_�6��+�ʢٿ����a�� *@տ��P2��{�;���6�J��?q.�q5\�3��C����چ���x�[NC�&��Q�LwR�5�k?؊K~�KM�T�X�3,4��A���9��~dCmO��"Q��������_jn$�;�!�#��sVU�f�a�Y�6�����@�W~3� �h�_s0�̙�\�1J�$is9h<�D�A͔��T$�z��f�"!?c�х>s'U`����q����.�56�g�J"�,���r#�~�g����Y�L���H+"�z.���ưX@M��wЯ�3&̡Ph�j�h�3��>{�~�R��w`*�e֐�jƶz/p��ϝ�|u��|N������������	�'q�u��I~�(��1`jg��p
�p\�u:z6YI�ｭY?�b��T��ӊy`L����'l�}8�=dK�0��{��R��O�$�y%�"�e�q��gCs<2��W�7��(�FT=<�����%��d�CY�>�P���5ڈ�qCIb���̭��k�D�װ���YkG_SW��h�^q��:��C�w��4V�y����&��_JL#y�ߛ ±u2L��鹏{,��ya)6AQ�Ņ�0M ��E�y�e190�Қ�[p�5��;Ϝ�l�h�YC�3����25)��ǯ�I
�S�R���m��7���}�B@�%~8k��9�F]�2�(�񞷿g��TKI��������?q�O~�~��}mhT����zSE�XEO}t-i�זA��q@�q��NRvk�ɀ��J	aIq�''�t�j�����L�W<w��-j0��)d�x��KOh�V'x��=�����z�����>w�5o�0O��&$)ķ�mB�2l��p�)~ �"1+���ra��}�y�F�ީ1�H�9���i&�^�~(� �b',�8\��^��Cp޹����� ����]�;L��߉+���"��3�ߠ�#Ҹ��9|�Kq�MېESS����-!7jaӚ
^�����W��֥4�ַY	�6�
��p�O��7.�ر���F�}�����\�}hm�{�F;h?��_�l��G��s`��߂x��
]���X5����</x��X]��.��fq��a��}hsn+�ЋE�Y�6,�X�a�\�>�K-vu��TJ)7&�s!�S_�.PӔ���`"^���=+�� �V�Z-�E2�Dm��LS.YJv	L˩e�y��x��Nĺ)�����aǎY���W���~��0��(�
����Z�� փ~,��iFH�!���VR��lF�B2�ߒtK�`�8Cp���XV S4�����v@�:�n�u���Rn^̦Qʥp�G?�OT`�L�nf�*�Bl�\���q��%�z \D��
ax�}7�����lv���8*aQ�7��jcv~K��C1X*��"���O����â{8��<-@�Qg��7͊c/g�Ry��g�p/�;�`qОC.�ǚ�S8��cp����'���\yġ(��sfƓv2�H��p�����l����쩶��� �tʶ��{њ_�T��5kעę\���Z��k�ɸ�ٔY�t�.�X(�Դ^�0m��r/�Y%sL�,�CV[��TM��k��tzh�/ �h��}%�W��Qm���2�4N4YJ���uUt(#��q�ږ�qz�O��8��	¼�'���?~�v����wőO���S�Y��e�	����|�\���@z�^O^�,2X�k�@�f!�T��+$�IO��%咼��Ixx-Zxj%�m~�2D~�R�����(pa��#R���^��f��0z�Մ���&n�ڳ$&SZQ�>rcDn����>�65{R +X��(.���м�}6�l��@n��(�P��z��f���ƹD�8�s&(�z�jcB2c�1���u��Ӹ�X��&�IX�!VD걘hq���5�l��7�a<��1Fn� i���S���6����c�Qaɽ��\���\D���zM�4'���Un���G���L�,�T�6=s�7Uג�t��0^��f2����c ���2��=�X�+ �F�}��슑�@~sdYf�Aa���?�0|��gb�%n����z�)�3���1Ǝ�p�{����[H�7!͙ř��a�Ɖ�9��V����~���}V�QR��CU&��;(l��]��fɹ	!�ʒ��8��h��Ұ/G��	Hؗ|���tyԡ�n�;�B|���bc�"�V&-X)����K��*y���m�j5���~o�=�C[��dM�_qA�A�c�3�1X�ջ�'�L!G�]�"����g����ͽGþᰇ�O��{��2�����֢jeJ^�%�Ϣá�ή;F|g����P�v�S�Xf��e�������ɜ�٫�Iu�{�uq�#�q��m��'P��ʗ�}PG�����>�To��k�¡
i��J�>��߻Bb�J�C6��(���a�*'t|DZ����:����3Bi�DpJ��n9>JF�0ϡ�T1/��zɠ�I5{S�if�Nϓ4R}�P�:tj���֫>+���-+8�Ҭ�ǟ��g�Ay���G#�k�	��;��p�E��̠�	����o�y�~56���Rm�^O�1m�L۸�ۗ�*��2�;n���ޅg�I{)ܾm�����m�S��=��5<��C��׿�;�)XU�B�='I���{�g�2.�;�]�ŗ\����Ժ�J�D��9<2oP\��[��\�	t��g>���Y�$80���7����5utM�Zز��s��ex���앻�V�c�c�c��=h�{"�d���"3SSX�v�4^�������]����A_) /��8�bxd-JkK�a�Wap�:��J+ղ�S'����N��j}В�h�Qg^��zu�Gul�I�'��rVMeQ��ĭ�܉��-����e9���krz?�~��yޭA�{גy]���*a�G�,��g�	��Mb���-�Ќ[�'�=^�\��1@�dGyPKX�䈕��,q���LW��7��Z���ê53(U�Z�A������M����n���Y�:e�p�����%ϼ9����=nX5=���> If�簰��珦2ȗ8�1�LAYzRJ\ɴ�ywi��Uɼ?_�-�122�7���YQ��vc�=����a`aR�%�S-T'
X�j��	g��,��U/�a[6�@ɨ�6������6��+��϶>��QES���l32��Ѵ:X����J�V�AQ���sw�l6D��&>2�+�E>K�@��"�J�0JyS�ʫg��f�iZ�֔�!d�I
�>�πiwaр�HO�/У	�eغ����q�{l�����%�Ϸ�o =jb"���O;����"���!~�=�^O;�T��G	��s]�_<���K4�e���@aY���4�>�rm��	��ZI3 �hB�։"�U�e���oF�2�0�y1Gc�7&�U�E=�@�8���:c�7T\�5qK�o�X&q�*��Tڭk����i���0{y�i�XV�~1Ⓗ�u�qE|$�����
[�;e	w0���2�Ay5��#Xg2W7óqbh}\����ˍ�,Y�p>/Z]Ѥ(q�rs1+���\&/�m�5�wK�Y����s�ԝ�,Х�|*�6���g�uHd�^̋��?l�MΎ�.u�V��v?$�3����i1�I� q����J���'Jr���V�@�^��f�������h����6t�P�����>������Dh��U�H�=�+�*՘D`Z[�o�]�<��g����t���a�L���j߹��q�3R���}�^D�+�n����VO�/��kY
�����i,O���&�/\����L*>JL�,8HV|[Gar���خ1_���]9Ea�%�ZB߽ǎ�0��4�?򜭠�_�����q�9����]� SroeY�"�W���=��䭭>�bu���(Y�)o4��T�7���$�
�:���o?��~��1���B����L��]��� �N_ͷC�P�z�G����+�j]�'�/}�Z�j�v�K��w�[a�M�&}�zNʓ���y���BD���1�Mw�%kJ�w�|岀HUq�g[�r}���Z��)H��G�r�)�e��-��ӷD��l�*��ɜ�Z���K,^�yI�$����I&T4�jtimi�jYb!��q|S��Ba��R�S�7J���e�d�=������Ll�$�t���;ߵq1w<��W.�?��7X�-����S��:n�l9&��ݷ�/|�R\���Q��Pʧ1UJ��c�{��:<���Paa��ݚ�B��,bMǹ�x����.����)��f+����)�j�Op�S��^D6E�t�|�i���`�����q����܈�����2������L���l�6O<[�tՑڦ'�e}�E��b����[��W��ѥY���
N�D�*��1��W���u��9	�rI�LZ�6�ڭz��I'[���5���[��6��G��2ʙ�H&˜U�G}y	�v�6��Qȗd��;�z�-��͏��E�+Ib4�Kr9�׭�S�>�2��^ȶ�(<V��Z$7���nB�d��UIeǥ7���|h<�[M��qк58�����C�̚52�=Ha��\���ǣOt��T�α�����O)���^�{Ef�E:�	K#3(����`B����ZM��7�D��,S��d�9���?ۡ�sCYSS2�{�c�,h�0Ͳ���B�>��GQh/��6��bf��u�f�n�Z�_�
��	�VO#/�jf$�2�k*�}p����w=�fz������}ٟ�L�N��(�]�d���իQ(%����`��2M
Zxos,N����Q��^��]yK��������p$μ�"��-q�U�/��t~�fKzL�O����d�G	x�%�!����	4�B�� �|������Q��S���:�yc���!���܇r�MU���Q�[��Y�_�	��H�d���[�%a]�g��s%=/"%��1�tdƴ�#���(�g����́2K^�i�e%>�O�D��@:N,�~����$f�C����q��k�T�q�!�l.�*m�#O���4K�!s�EP����\H��tc�(1��� � y�3�d�.	o��>&�|���SzC��-d�%L�Yזtk�� ������*�pO��{lL�'b*&<�ޣ�d�fqZ��?�J���l�9S�S%�\+_�]2u]ۏj��=^
jV�����-�qJQ�@br4�)^3�Yd{EW�~<���1`*vb�u(�cA��.�d){uT�s���|'=�(�
W����8�H� ��M��}bL��%���_B?��|�|ALM4��q�֭��|ƍ��
��/K���h^�����������o�	{+z=��1�쬓J��"�]1�Ë����h���X�z�f��|�B1m�b��G�/`/_g,��LP0$��S�sp"#�ok�����集"qrGC����b���n��Z��⊔�
A� NR$�s���}�ף�&��n���#Е�2�E�6��|�-x�Q�(��5�IYWSp{EWq'K%�$�+�;-)�5��+���3��tZ|1���n|�{�c�CC$-�n^��l�2���IE���<M'F�G;<W9!J.q�e.^�{:w�ꍼ��Iq(�0�L��q�gZ��b�Ԧa'{pJ	YKȘ��_�>�Y��:�D�R߃�Q��u�'��Z-��u�ku1[W�|N�)�dy��.R	��M�s�)G�q�]V$�m�I�{�{H�����
L�}֗T��^��e�90�s{��Ǹ��ߊ������{�,aL5	���}��W.�oo��t3��~������9�l#"�)�U��t�d)P�#����0S��_�*�ķ��iFEA��Bʸ�YBj��Qg�z�8��g��otm |�7��߈ٚ�����Z����8㩫B?���ĉR���C3���������[���o�r��E�JߦU���Ç˛������(ɜS�W��-�P��@�T��-lP�%s*��t
���P�4������r��r���p�^��>;��kS�W`J#I�K���b�f3c}N�U�����	zr�'���5��y���F#ڟ�?0�DU��~�`E96:��|4��������2�ߧ����G��B�Q�����W�2�A��^��&JXV���U;�<e�=������rxz�ϺZ��+3ǡ cE�F�(���5B�.����c`��J�?F�N��5%0�ڢa�F��\����;+����}�lY[³�ހS������t9�[12�N`� /2�,R��B�W���|�G���;�h���э���g��T
eLӝ�ј����$�֮E��@����GLF�J5�r�����z�KKr�V���d�t
޻!����p�'_#G����Q����H���򚉙����dƂ�x�2���7l���8ë�~g������s^��U����Q����{�o\(}�/~��qʉGa�:)�����\�?<ZC�PE�\���Uf�R�j�"镑�6�3^ љ�������mq��"�49ݕ}�a0�����Ey?sUd����$k�+��I�콆����^`��n���N����k��Zx�Ϩ���zk�i�����$7}J	���ҽ�1��	8��?ƴ�tD��-5�do���ɡ\���t	����s�4y���]M�&qe<��1�c��`���k�blY`��s%�K�#'��~KK���;��M���#E]�� 'I�SOO�T��D�+IL�b�NK��Bט��۾�4~V>+}^�.��M� �K�}K.a3��'�`���f5�cq��x]���b����<.��3x�ZM�8�+1��"���Q�$����(�p��v�ß����1��-�tD��e�Q�b�x��wF?�@P��xĚ'�:��L�^ºԍksMW�8�O2*L�3Kky�^��z������i����B��X�C��'06o�
�-ə�ar�K_3|�õ�����E+�,�T�Թ��c�}C�HG�~g}��`�s+wI�C"��N^�3�{�{`��JeZ�Y�h�V��Q�/=�Go��~6�{�$�,,�$_���6b$S��$�K}�IC�`%eo{�_Sӱ���,�^s���k�`o-�8��T��Az��Az\X�Xkj#���3�N���A_�Ƅ��s91B"�I�n�:��k�Z���a��%��Q
���j�So`@o~~�l+��"M�rb���8T�I^l�?^��.�a�u:�ߴ^è�12=)�'9��"̝Μ�s�z:5E���1%0�v��ot��0I`��'�c�z%�q�=��`�Ӂ�=;���7(���G������Y'l�5�7��8����qۭ���x�!��9g�%���<��d��%r8DmY[�\�HbӢ5���ů\�_��~,����H��GV���`������|�0\
dL�����.�B���SO܂���M8��d���P~.mD�c��]�{�c��|���qѥ[�N"W��э.b.>O5��9"e)�    IDAT~^a�B�!�lq���@��&�&�#-��r��8�O��������yzȤz������8��_��rZf�5j˸�������°�8˔^��f bA.N��Jr�|h�0.$����?V�JL',f�'����(1]Y�����@�z}D����7V��$�#z��vD�#]�M��#a�z�Z�'��+O��Oc�b{�Әk��O�0��;V���̳��=@��'Л��@�T��ZC{�9�7�����/.�60�AJ��S(U�(V+Ȳ:��ɚi�hs��P����&�KR�L��N��2*�N{��8�5��1��2>Iy���{�VGv�R�?`�h���� 0�M�Ƈ�q�w����It%�k������}t'j�s��T1�a=r�2�e���� �Uh��t ��z��E)ް�"[-���D�LZ]y���j� ��}����V��%�ސ��M ������@w9[b
�@�c_!E�T|�k�a1젔ia*�����8�eϑ~p���I���~|��X�7���#��If��F��n܋��O�خ��
��?�N�iy�&���������t3&0�P���&��r��Nl�(M�������6�X�<�H��ґ,�b��ج�Z@��ܑ�z��
����;C�`��i\��4��,��-�C����������TcӦ���5X1e��=�(��ן����Fr^�Z�:bBC��+��y�lIaT���l��i�2���pbq�ghR��4�0I�~���/��?o�O��J���H�p�
$C!��f�~�DU���]w.Ж�E��x-��c`ke���+/oKwg����B�+�O�Ǩ���p.��gp�ZM�(��B�yxA�o�	��>���B+���Y|�s�A/���#c*ɤ�ta0-3��a���i����"�'*��uE��\�>�����Y�L�<vC����=���ԨJ;�������F]�5f�ݡpų3znWm}'F��EK�J�^�hc�9���醾��`��3��8'k?�;�'y=��9�veE�-���o��9�0۫&�����	Fl��s�=�Ͻ6d�Ful���S��S�qܔ��J�S�i^cw�3�C�b��F<fX��{�c��$�'�[ _��V|���0*�E�]Y�b�`�X�[Le/�@� ����za�c�c~Ё�&�ۧ�Ed+�8v2묩Q�c��[��0��9������ۨ��lZ���Y�eMq����iQ�q���%n�Z�(���"��WH7Z4b�$c?S#�&&���"��ȕ\#���o^4<�Y�����@`:�"?�:Zƫ�u8>z�+������}|�?�W��zO9j>�����o���q,���>���ĝ�߃���s�>:�ش&/ɭ���
qe�\��$H%�'*���7l݅/|������f�������5`��To/����#�<�E�����_�{�݂�%�֯�ģ7�C�~#^x�Zu���M<�� ��jzT�yTJ�i����� .�эX��v{}�LC{g]N����Q��'���Y�*8-���LR��i5Ne�:狁��x0袐�8���l���s<�>t�+��|�[n�_���en�(e�����V�b��J��{_�Kn �t��plٳ��xRu�2I�쭐�1Qd�/	�/��jG�.#�9����E kI�i�Gf���N9�y�8x�fT89�G�?��s-���>\s�}رo�6
�X��M�2��J�=Qb`J/��ի������%�!_ʀMJC��� =�TL�Y�`�%� �J��	�%��aW�Lɘ��e�C�a�rM	�F`�X����/8�8��Xo�L�����&��F�_n�s���x�q왫��M��*co?��A�|�l#饵1XC��k�0���܋��됛� U6;r�B��2�A@IU�����/���}���VM!3QA����gL��K3q�폐�Л_��/r�$���T��j�	I�Hò7V^�/}�I�Z"��!4p|V�Q�'S8�U��^�\L�pp�aY�|xP�-�����f͌����n ��6|�{�a��FjH�}Y!�B%�5��C�DrkYOV�}#ɓ������М	1 'RsJ�-��D�ׯjKtd����B�XY�����v{��F1�kL�؄�y�O���(�:k@���&�>MJ�Kv4�z�,VDq+NC�*��\�Mv����֗R��)0�JP�Lj�B�9��;U=p�P�d<��Һq6?d��v��G�j�|F�>�ą� ���֥룃�SŸx�;�ٷ��0k���P��EJ�>ۓ1��s$��'��S��>�3��I����V��*�����m��]K�z��G�9��G���xD�f*dGT.��L�v"0��?�8�(s`����c�V$��kK���ϟ=���?~�aq����8Y�����n����Cv�x� ���1��I�y���r�����1�+��{K�
�Ƙ�EɄ�6����*������Zk�� �q�a���T/c�H�$�Jz�u�M��������l�o���h�(�Q�t\�")իg��-V�9-k��a�gr�#L��X������y���-�2dG-T3u��ͯ�˟}0V!���v ?���s"~BI/jH�=������:p�#-|��˱m�2��5�T`�
ݫ�h��U�u{��R������lzow��-��=��.[�()f�g{=6JT��T��F-�#M&d0T�[���4n�7t��O��ԞS��,U}E����µ��C���"~�_h�dDͰ�!Md�Tv���@�rT�m��|M�|�I�pÀJ799��GmL�x����_����vF�Q{�ƶ��8��Kp��7`qy��������m��Ȧ�k��Ǘ����&���O�%�|��(�;k�vO({�ޜ?hbf-9�"�]��k�߆Π�F��'ώ�������oz����Gњ|L��+���[1�<��Ԩ�'m�ƛ^�'8��#1S����G5���C���N�_B�Ւ͵n�jlܰ�v���LLW1� ~z����U�b��B�2�no��)��"�Zd~��\��TiM�R�P��Ê�3{M+ժ0���3i�-.�yOd���ʍ�X]��O_���3ƴ�Ū#[;w��|᫸o�v�Ry�cF�^�+xP��C_|�Y�*H$�2�R�|x�W�b�R�ϕ�N|��LV&�uyϨR�KL�L~&3�q�Y �}W��Z���y��� ��b��g���&���>�+��Kݜ�G��ڍ=��%R�P`�v�LNL�������_�Yl\��A._PC%����}tz]韤ĸ2=�r�"��r��rM�RQ�ى"�d�� v�d]{趖�,�5/<	�|��XM�.���/C�X�8��~�C�������݋�w�W1(� 30��0T֯G���@�{�'`6�	0�4�Xع�{gQ�VP]�٩
��,Yc�B���#��'�t�����a�mv����$XI��Qw�ɾ0��e�P�!O9o����0�9k7�j��}"Sh�[7ӑ��$�'��bNz�Ϻ4߷'@U�A�Q��r�6F���J�ox����QJ%V��b�MXd��=5|���7lC��Ũ;D�iw�"�a��ՓL�\R��<8�+T�p.,硚y�I��@�\O�F�>��H�I��OFl�k5	��"�:�T�(sJ�9��"��i��cɫ��(���-2ڱ{#)|��Z2�Y���LW���*��^P)��i2��S���&�	��]b���0D@)�>L���缒���ȧdK���x���ep��?K\s`3	���y��?���%{��17r-b������9��}��}�5�/�z����`�y?�'�*��,���������n�����Q�ŃI�3�-!c��*ݏ����ف�Hv k/�H�W�^v�Rl��Rr-��H<����Q�"�|�Q���Ĵ'1�fb&{DJ�&_Դ��,��!���-~���ˮF�J�T��YY� �<�C����I">���8�R�l�߽ "��d���M���d�|5gL�]��"��8TIz��YL��)�Û�@�t��>�M�|?��"��YB�����r`Lm_���N�4�5bR���'��q	{w�m|�$�H�z����
�j%�y���D./����{T®�d�)3��	C��E��Trn�Ơ9��7M�#�"VMVP�F�P��	x�e�& �s�G*ٟ��	���K��빡k3���s�F���z��>ڽ�G���U�ʔ��d*�B� Q!�C�b�W�|C�*Z7f`)���[�H[J���x������rM!Ccˉ
����z��k˞2ﷂ<5�fr�rr<Oo�~�%�i��T�`�0�FKu�d��+�[W��`��SZl{J	k�٩=Rvڒ?�&�7V
��2�$��̋�	[�x��t�>��=%�A��e��9G�c�kT�;u�����8��K�.-(0��������S���6|������3�݂/����Q�LHr���H�!�\�A��WĒ���Y~C��7���<��fg�N�E7dd3��8��/���*����o���5��w���I��j�P�q��qĖ5(������ݻ�s��-�L�+L��*_(arz�֭��u��K��}�v�u0ʖ��P���Zu��t�
�A�U���D�����F#ȠL��7��.���5�5{�]l�N��~��F1I��G	���y\p��p�m�!�-�hnIJ�GA�xv��МB�gh�[�<-����X�����5?1�O���v��L�QW���*l��� D���������	5̓^O�ƍ�����O=�()�(�/'�rF��~�]q{e�(��ܴ��-6�j����4+�����5�1����>旖�g�^�{6wTz�$���l(??������6e��*S��r.0�߽�Ӗ�bR�*Σ,f�&�`���P
�,����z��8��)e�./�D�$��L�t�������o��wΡ3,�7,aP�Vo��'����,��s��dMy`�;(����c���h�ΣT1`:]E���Y.5t�0#�C����Kh�����i�"z|�t��#�z,Jd��K��PS��-��(JM�D�+�8VX3�O|���2v+�8��	5�/��k>�^w��ՑIu��-#5l�M3x����iO?
�EGq߆LW��Mw��+߿��� �:#�4�p�W�L�qw�Q@6,q�ԱAtu�3s������DU��h�pfH��i�E��� ��e��1�ЭO��%���5L��P-��������9g9Ԝ�ԕ)TgVˌ^�Sw�uc��F�Kll��V�qk��z��\���L�S�g���X���$2��S��Ϋg�^ɦ�Ul�K��k261T�����0����x�%"�i�@�L
*=OZH�!��W��e	�ފh|M�
Qڦ�� �}p��c?�ޙe����R�w�eɾ�h�a�x.H���x�L,��>��aS'Q�w\�좄��)3��f��"� �s!=�;�s%�xvi!��a�g���r������g��K�}�,�� �;	�*7��F��/������;x`WmT1Ls�ؽ��F�K�aK���V�ґg�,}�0�gs�x}IN�a��G��<���p��Ɋ�s�Tů�R{#S����I�E�Um�H�˳������s�e/�;y�Q��Y��Ud̗��蠿t3*�0��L�}?ŻB�K����=��^��}�=��{1���Z�5Iyr|H�<��x���F}s@���^c�Q_�[����M���J��kRTY�g���1�#� �I��9���üN9���b(Ag�f�Ȕ�P�X�T�����6W�1u��oA����2������>B��.~���Gx���Z�*�f}�G���E[Y��jχW+y%2�Q�1jwd�L��@��R�%�2���)aXȊl��O�=�^�mVd�)L���j�K�;�AefZ�.q�y���y�8A�)[�Ș���jD���1ͣ/��5�y2>���bm>)�G�%9]�����4��_��U��e�����=� ��y�ũ2�Tͅ���.|�����܋׽����}k�@�+j>�,�=�;% S(�ň=���=���/����6P�y��4M}����?{��Η����j\��;PkjŦ�m	��j��j�7��^��ZmK���w��:�7��8)_(cbr��$F�)th���D��&6�DT��ϡl�Wє�a�O��"m`Udv0�ZS,���H��`2-I�V�������uL��5�.�~���g�i�7�_|w��.��ضm;R�8�j���s���s��%_��9�U��0�J�~� 		A^����5ӎ��*���z��j]bD����IS8T-0�9��6kZw#����.��ܓ��1i"Ì�'\�������]�2�,l^��jt�\n��� +�H�$0]=3���i	��V{��ʜ'����g��逖�K^��B��`��6�Mw�l�SҗLC0�fM{LG�'G�>-V�ϔ����F�
}<��-x�+��#6P�A$��gR�\x��g�����?��m�b�����)̎�H�:�l}�%0I)�h�x�w����?�8�s�(W�(�[��L�b])����i��ʘ�D�.�5�(�k�L�灌�R��Q_L�h�.���
�� �9���%#� ��U�lY����Z�`[$���ʽJYd?SfI�8��h�D�� q'�ꡜ��#��SO�s��T��a��#����J��{w⒫~�_�p/�k4�裔N�B�v,�}������6�qm��[�O"��dUy���4�Nrd0�������r"3�aHv:�k#�m�4h!+F-����K���TV
=�Q_��49s������Gz��3a	�`;dl�ɑ�l�kAj� 8{"̋�'7us�#+�ɱ$.��9[!N�:�.��2���W�d�
�5�k��&�Z��P����15��_a'�T�U�ʏ��G=��,VG&L�d_���wQ��᠛�D甧�z{b�������g��b�A;��s;���4�g��)�X}O=����e�1���@�+/t���B�J #���T�`6Ċ4�:0Uz��ʕ��0����{lL�)0��L�﷐5����sN<��W��'M�d�Bb�3W&\ڟlds<�p���~��)�Y��Ō�.����L��H��xW���w�j���T3����|���g5��S�9@��5g���\[�Z�3z��^�
�!@W�R�D��Ÿ�a��K9}��]����*w�v3D���X���yϻ�sۿ�+��</�x��_�U�%�3F�{���
������y�1������9|�<�u+�K���8��^WX5��
���G�� �V�^�,��+ �h5�#��ʖ�/��$�{��` W� ,Pg8�����'e�.'�sT���j�EB0E�g�a��_#ULU
bg�����h,�#��6�w{<�2�2Rż�zEOa�-�����g����"? �z]����u�9��{�ǀ�E�,��͉����<�|f4�̍2�՛p�C��N�)�KyrJ � �� ����I{L�G��=�����T�}�]��%c��?L{#��R�]���k��]�}��8�ȃ�7�y�F������6|���ే�����IlS&��2 N;ƃ��J��!� �&��:p�7~���:�F�|�JiG\E	L�Ϋq�[_$I&_�������⒟܆Z�}Xگ�I��nU	O�4��
��:��nW=&�\b�v=:6rto*����Z��L��*La���I�%k7L�dc�ٵor��4�k�*.���)�Emv�2�U292BD%;�[��
g5QHu��/��#��S�Ɩ�f0U!{����~}�opۭwa�K#���pA*Hi��.�٪<�v�N8zQO�U��1,9���k�$���]�́h�Xyu0�3��d�D�6��3�j��i�y�2 Z�rXeT=4����<gd��    IDAT��*qġ(���bO�R��ew���GmXF�P-��"樦�5��i���&��P��151�
��)4�Y�]�l))�s���M,-7�dő~8@���kjf��r���];Θ*�9��)2�^��T�Ѓ&p��㈍�8t�j�q&�[��BY_͕�HP�/����[5��1���؇_߻-t�-L�τ?Ci��r�����a�ѝh�/�R�@a�jdWM`PL�Oc�Q��h|��ϔ᎐nw1�_Bs~#���Ȓ5`�S`:`  \��"�!k
V��H�z��-"�b8��=J��o@�{������V�A��?�R�a�`�w�K��<6����OZ�C6���=O�Qoca�f&V���0���c�9�u0j�.��f\~��ص�!��'��>��N�\���׶5Ie�,��l&��539S�����-����㿻�.+Tg�������)U)�@$8h-���Ùg��5:�G�f���(��Y���X�����Gس����م�n�ؚ/OJE�Y^-N�~C̭J%��52`,�)B��4 Y�0��M�\�D�|��b� �u)�3V�D̪r<�L�DB�$�V��$�w $@ۿ;�z�+�K�1z���}�c��=O���L`#�ت�n��+_7��$���/iէ�����D:J��SH��h-Of]�����1�x���C������t.��Y�3Vb�K��sp� _����g"0���K���΄�N�S���/V�v�eJ���&���Fi�(��'O;<�ز.+EC����U7&��j��>���^s+��2�����ʈL��&^��x+���s�1%����dLO i�yA)RKioe��[�r����,ӟU��xⱇ#1|_X1�_����
��#)T�S*3�yGy�B���_s�@��9��������s+)��}qp�lUR�JrcJ���}ձ*���H�^,Lڿ��r�'���
3�7�x�'?�{������=���b�K,ܸ��Cb�?��Tq���Pc�!�7]�z]UD���햀R����s8��Ux��a���KEt{Q]}�-h����(W&� �J���+-#���j6���9�@��;����u��V��3���D1����Å\ۢH�7�<9c��z$Lf!�l��.���Wё��+���>�aeb��d�;M��u�� ���l�2�e�+%���Fe�,�kڐF!�CZ]t�k��a��i�*e���9-�90U%���`�A�R^�1�0}�iG������B_�� )���dL��E?T`z�����ރg��)�?ߊ/~�"�|�a|��oǟ��(�><9q�9�����8�� I�H |�e����b�Q���dr���E|�����B�pΔ�����?�G�`��CdFw�F��M/Ó]'��)�*J��P��G.,�L�ɐ�b_�r����������;�R�f���ce&��H~B�ă��g	�Bc��Q�%��+sƊ&�J�{Y&�^}#��oa�kbح!?�cMi�M3%��ȡ�K	�n��X��G��Ĩ�F.ǹ���fQ‧s75��8.�*@�Y��M�h[�E���DhUI���ʦ�*�I���]����{ۣ�xAS�y�Cȃj`O�Q���r�A��U�U�x�18�i'㨧�re�T��;����5[H���`��u�\Fz��oh��h՚2���#��L:��/�s����R-� jvL�ut�2F�vsK�_���0�D�� ��bzՌ��4��|�n�#�ԝy��i8���dS�
E^�w���!�[ƺ��lX�-�����q���X�z33eT9�rn�������o^y~y�.,��豟9_0s0�3`�PD����Gv���R�	��� �j�R��:�r���GJi~�����?��]u9l�P0`:!=���H��DΫ�2���T>gL��H5[ʘf��T
C�V��f}��fL�)&&,v9$s�'�yE��ƺu���X39�8����Z8���q饿�U?�^V��Gn�;��:���'��o��1\v�p���SO<^�R��REIG�FcI�H,ש���[ild�5 v�����}W�t�BEd�dӕU�����-��x�_�7��Li��C�@�$l��<l(����y ��[�����/�_�]�}d�3AV��a2�F��1�� "�Rd����祖��o��P�����i�acn�f��#o���qQ-.�INج���d&��z�f�/���c��|1��q{e}�0Y�P�Y�i�3%�<�	�;Yg+���X�"�@FN�rE�F�l	6��V ��s���%�$l"�3*Lg����^�8{KaʜDm�^س��	=�V���ol�n�ki���]�o�5`*
":Z�9����w�L��U���k"�Ow������?�{�YX?����{"���E�������7c�vYY]�n�_�^:E���Q��X~��%�AMb��D��(E�
��R�

Ri�L��w{����9�����<23����s�w�{��ڗ߄[�~��H�!���?+2z�"B�a��f�Hw?[�9�߇���e�8���G	|ܛ��F���1�2�(���?�*��9��wIZ��H!��K�̚�xe�P�N��Cy����P�Ml��a��(�GЙ[�����=����=�һfy��ΘF�r��[���z\��!H_��ɮ;�>&q��(�u�3���rȀ�(��:\!�F��V�E*��b�ˈ�I�|V��N��O4�,�Ļ��r���(�80��~�P�����l��_&+�=�Yd[��(ڴń}�.C�v'������Q�Z��_\=԰���3��U���+�n�5���s	�+����LJ]z�n��P2��0�V��١)��	�YjK��j����g��4�A6�H��QU%#Yģ̚��m	dɘ&��ԛ�T(�m���ǐ)����9-��
�<bC�)��sK6|�A����`�|�A��[O����L{���]���q�e7`fn����w�YO�(����W]s;�����k�6|�oߋ׽��j�b��.j�eb�"�pHF�7�R�L$� ��_?��~�k��sh��H�
��&�����^�Ɣ�0�9��W���A���9�� �j���G��JlX������I�����v��༯^�{����	kE��r5���d+���-��7f�a��+���!�a���Ӫ�&���0�lb���x!)�H�l�w!�G�����d`����?�*.g��#v���2�q��=Km"ָ��U�<0Ƹ7��Hr��Vm�C>��şoa6:��
Otӥ��Qv ���g���+��/��zm�v�{�lG�&1�l��������9��	t))�H��kiZED������5��A��9��1>:�l&��@������v153'li��U�!q�e�5MȘ�I�){�	L�di�m��]1@��W��G)���D�l
�cE��-4�s���,N=!��2}6���jr�&ưi�*�p����?��N��1("�����'��W�?�m1��NSALڃ8^(0};�Q�؛�+��A/�D7�ɤ:7Ea�����L�-q�%�ʀ����(����R覀FWG���8��W��ȁ��.L���2�&�d2 �������N}M�Z#.@�4M� �4"H��b�M4�O�է�����|��0�ty�	|�һ���6vO�`��"�u��x��'�5��Ԟ&v����k�b2�,�V�?"`4 r .)ZL��o�9 �[��?�e�����e2�WS+4�@&^��~<�������J��$�(���l�'��wb,�aƑc�>|�K��^� =&�TU�̊���K�x��n�E�[��D��c�"V�Q�h*�aq,62�\�$6����^�\2�3T�d ��0)Ԅ&>���V�-_�����[��i�bsl (�p(1���48��k2p�P�� T["�s���E��}C���l�{ԋ'�����9�K��p"���j�ʌ��5��n("P�C�O��� �u����7�;�,�'[�|/��M��H?�?CM`�̋;���"e�gG��{�Z��ˊ���c��DSծ�׮�S�A�[�����y<�ñq��*�o�;x��=�^�У��s��d~}��K�ϏK��%EE�I���9���X]c��|u力�{%��g�j�H�ܶn�b�qq�6o�Df�C����`ҁe 1Ȳ@cE ��u*kǟc�Z}��(6�ܢ�c���x�a{}Xv�c�`?9������:k�=ቧ�x]�cieC�~�-�����(%��Q�7a
~X;(���Rqy�KsC&VB���	�h{=(V�_FW<z������K_]lY��C�)�m6�H:�t�y]�kqئ���[��	����']�	��8�(�Ĝ�z'�zN6``���CS��	�,a����-l�eB��4-d�h������z>��µ�F��w��O-P���oI�z�y��O���VM�����1�R*�R:�<	�N�Z��y4j�#K�ǌL/��R�Ψ�Z�e�{g>��yzK4�27�c�ڵ�\catD�A6-� ~��S���9�N�r�Ň.��6��ʃ�ꔃ�w��;�]zf��q��q�G��IGm�C�=W��v������$��S�/=E�SR�W6��h�Ǉ�/��-0�Q�E��Y����\%!3*]o �\�G�s&^��g0�OՀ�⥸�mXlfDi�NuQ�tp�	��7���K
0�
���������a<�輺�|��p�/�q1���)��0	��TR�CO�VNpZ`+j�{6u����<��5�<g(aŧ�Bj�A>�E����8�i�+�M�Ǳ���i<��v<����j�?��gY�ɋ�!�} ����[�G�E���pp���V�5�1ل1�^]
CwR��$� �m� ��K$��L\����j�Mdŭ�;RJ�Y�zmT+s(���g����D&[׶?�i;�:�J����*$JH�HP�+�r��U�n���GG�L�Z�y���Tdsi���
�2�������k���G�FWb5JI�Ο�"���qaL�L��4+���=��fpap��c���>��4�'�"	o��1��q���&ny��������Ux�+_��?�Dr�<����M"}G;�����[����`����(��x��T���[���g9�P�^)���K��QP2��k�z`����%D;L`ښ'�0)���)�2�-ޣ��[I�XM�Q'Iq�M��h��	­�Tl������q=E2-���:���L�7��k�.�2*���|z�?�8�CP�fBؔ��_��j|�k�bq���d/{�I��G߂�+x���=��vA-x+�Dk��Ag�@��Ǯ�>�ٯ������E�8�[���F�a�=z$ ݫb��,>�q[ǭE�]c�ʁ���[j���w��>�B	<2|�?�m�݁~rL�e�ș�L� ��aI�yɻ�ي&��J ��(�'��N;�# �,�$Б��7_�fՙ�@�0��Q`�]cY�Xg�G��_֒��5h���%=~��7B7� :: ���r�(q��1��j�2�5�k Ә���?�b��Wس�=�Ɍ��/1C�@'p-5�W��`歬]�*WwN����0w���o*Oɪ;z9����Hט��v&�=�cǛx��D�z}�X���UQ�Ӭ@�x1}����Ó���۪��^D_	�ɨ�4�O����!�C2���<mD��T9�?]���u���Z)�D Z�� ���4ߺD���.Y��\B�Q\���j��h��)$��N=�ĒH��y�/�X��q�2�������vhT6�^�v��P�����M��sv�z^Z��Z+�Dw�� 68��K�3�΋B�ѹ�HF��Mz�^H��}�R��"���z>G:yNb*3��̬��f]7�T��Q�=-/ʓ��n�z�N���=h��ؼ���^#���"0�g<�x��u(�N"S,
�h���PC49/�)2�S���ޤd�3�}�H꺂X"�sT�R�5�a��.֎�O���e2W)�k���HP'{�l�*�ɤD:���g�_j�,�39�RI��z��E,��i�M��1��vt3*�8IU��tr�^���F[�Ɠ1�6�r	L����� ��ƚZQJ���E�A��6�\�sLS�F���R��c�A)���ލ������,9p�����	O[/��.��-8�kbjד��?|�z�ȱ�a\5��;ԫFq��!����S"%K$�1���|�S�c�LG�yZ{%�$*���^�3_~�2�1S>�Kp���Qij�$��`�*�w9^�W����m&�-=��p��
(+��%�
6"�t��nَr�Y�KeI�8�^�#�&�$��yY�.��T���A�����Y=��e�7�Y"�^_@H:�E>�F�9�׾�x��YGbYY�Yh��x|�\rɏ��?�N�	�S:�i�ڢku#�x[�ӾBew�
���ś�5	2V��h\e]R���}��)0����WxPɽ�{��Rp��9��ܪ�R��5���tG#pt�n�01V��g��Ï8�bA�V;���݊��cl��Bv|:�"9J�HЬ(�A�����j�2� fD�D��c�� �@��f�dml�X�ӉW�:�� S�wJiG��l��p[�Z�dL[���^2�\>
L�nH��|1����T���tk'2X;�ź�(��(d3"(/�3)e�B�a�j�����4�������މ+nߎFf��Jy%�&@Dʛ��1��ITg��}��j9r�1��rR���L�<J���T�Nϣ�P�����Q�C���=�6�����|6&���i�5zhN�!�hE�b�=�\�u}����?�Vkr�.�� KV1��8�o9?L�S8։���4�L��O{N>by�qI���e?��ו��o�ƻ�<�C]��?�l�p�Fu���^ص��d�n��z@ı�GP�.�7�[�l����>�yl��D/YB"[D:�E�}֒��y&�)t��V�n<�7��4��G�H9����!*!.��{,�W��]w0d����y���]�[~�]�"_*�K���:k�I��9<^-��{����3��x<��W�B�s�wf|$?��Y������£ʜ�W�b	� � ��k̭g� e�D4�&fޢ�*�r-zx2�C�V<?{�ۇR��y,�� ,JF�B���8{�������~��#��Yr�5H��Sq��@w��'K����d����7��3�_�v6�6�l�q���H��ц�[AD[DLn��Z;T�z�t���
��2\����9ǃ\
t<���Z��fAU���O#I�Q�^�IS�U*}�&3�xL�~����{B%~������/�o����tA�ѳ:���֋���1���r�^�=bT������y���$b`;���C���74�	*�}�2�{����u+*s�5�c�̓#�7�X𲸤^ۗ�=��������[|_cx�"������=��iT�d�3E̹�>T-��g�=�37���̰��y���M�s '�5�yw&�z��f�&k~"��	O�o{6��Տ�nw	l������Ԁ�rL�Y�T���Gbo�1O�~)I/Lq��52s
����3�u/�U�����ʊ8S▶3���f��mAv?9:��GeN-�I�����-ڪ����� �L�Ţ�ʃf��9,���wc�ǽP�+Ƅ�|��zL�p>j�f[���9'�ђ�FG�"��N�۾�x�(P�n㰴�:���A�O)o���|��x�_ =�B� <�s��U����p�e�bna����w�#����k�]�|��ocj����� ���D!�F�z�kj��K�Ӓ�k�{�a���#&cz�=S8�3���|�j�\
�A�T�x��񚗝(�.��]5��x	~q�c�6Ӳs�$Z�YRML�:ظ���7��_��tv��ܛ��p�Ϳ�Ïn��7����xA�l��/��W/�{*)��ʞ�<�S9�Eg�UI��c��7�4���Y Si    IDATE��%Ʀç<esj�;ٰt�͢��l�~���#��LDSm�����gW�=-��~=��*���;݆D�s 	��)�w�Q����E5
���^_t�ك��	�ʎ�?�_-]7^��ÿ�%<|uK^�oZYH��8耍�ԧ>��	:�OJ�+�������_X�F2�D����/�H��d�.�̣]o��������}!�ܤ��0x�Bgo���${:S)C�L���3oY�yF��@��A�R�`�
���H'�����vk��/xN|�)lȎ�f�oC�������'�V�~����i�S�hpK�3j���w`���z�O�Bez^��i~�S�ʙ\V����ʛ RGgz��E)��}/S.0�r�|LU�_�@Oջh͐1�S�6���VSUmf�K��!���J=���2�̙yB�Zss�Ⱉ���5|��ލ���E�B۞����:~y�}X`���#)�O���7��|�+t�xP�r��k��m�=�-[���C��B�XF�4��;׌1�b����=����p�EW"]X�>g�Fd��x�4�"�e�۬#٭a"��чl��O;p����a���NY�h���}�ݾ��`A �I!O�~��9�X����oފ�`c�(�Kj
��JuݒP�F���P����L��7��o����1Z��"c�%�@d�9��16a�X��FT/�I��EH8N\<W�%&FV#�@��wI.-.G*�Cto��P��6��~�P��x���M�B{�&������9��(*\[��Z��S)W; 
��(�-$ẉ ���f��ٞgg]~mԞ��o���ya�fI1n�X.�7��KݼP=�l=IR�+�Ǳ`T��,|I/�#ot�3�suUB@��3��3터Ν�j�I1��ȝc�gEs����2�^����ܘ�[z�{�cc@  ��۟s�]�X���ԟY�D�+z"Z�r�娐��X\Bj������E�O�}��;և.��[|M�ɹ��� ��\,�C��s+̊D�P��8R���
�����P��_�B�?{�qm�����R+F�X�������D%(�rh�X��E�U�d���[���}&6o(J��oC)�����>�/��O�H�Vab�Z$8�]!��#C5Ib��K���=���[��M�kz����\��i/�����D��f]�g�4XI��X~H����3�X F�H����=�F�%��.߼��`�P���͖ ���9�)&0�a����;t8��b1��eȘ2#�	l��A���'�aK)�%����ڦ�¹*@�62�9!��i��@�?�׾�����ǲ�� L[������g��|�r\��[P�.긘����8.�7�B'�]q���ocz��s��qλ� �&%E6jO�m��x�������(��s#���O�ܿ^�F+�n�7��T��L��s?�p��'D���/����� S�|!�Fc^�5��;0���g��|�8r�:�z �|۝x�>���,[6�o��8�C�X�{���o߈��@�4&�+�2�O$�*o�E�a�� .�l<6)�vW�R(uC"	`C2��U�#���V9Ա���^|<N<r��}�Z��.����ߌހ��3��B�{n�@)��_�s���	�e�����I�M�r������6{��������@��O��/?t|M�%FAU�%�~�Q%�ߝL@_�)�m$=��z��'>��ɒ�2k�/)�|�F��ڻ��+���X��"tR�eh�9�6;��.�[o"5��F�Mt�!����'�ZQe�kR-�).�-��@)�4\���9̚tX�� �D��<�[ċN>x��0��"��3a���0�μ�Pi{��S]\���p��:���48։����8���t�����s
��Q�V����zi��j��;�$��\�J��Y������ˎ��cP̢��cʠ�Q;&ȑ�,�w��Ӿ��֛�'�5Q�H/ߩ(N8b^�D###X�r��C%+�k��ܹ�z��4�߼��؛q�JΉ틜���Sx˻�zh'�-����E���i�?����`���Rl��\�����a���㫸��{�~�F�E��-�<������yl� pLL��F��D'Q2e�FhA�����-�y�������׬����y9���y��T�$0:RD&˟�d��k��E/���5�lb��	�>�H��x��^�����d3�/_�\������	GҤ�f'�0��!&�6[�z�eǕ|~���I��W�*G��N{aȓ�X�u]�`� �ݛ�O)��I8�a�d�B�R����kOzt���*dLj�[S�p,�%�C\Q=Ҋ�U=���ZYd��C������3�аKM�bŎ���:�����1J�5Q��H�=�teS��G��J�@����F���?&����G%��ψ�3:�b2d��f��.R]K�=��OJ�Xm��_��T�Lb�����{��[!r�V0m��T�Ȃ�Sl�e�*`L�lw�>�Ҙ��������g6����~$0�����6^�g,5q�u�1��F*��/����� Y�>s3.��-f]��W��6:"3¼gXB԰��7�����I
nU������
@ѭ2���J�pĄ���R���|A��YQ���"�!�?�]t'a��BJL�#�ɠUo`~v��&�m���8�oހ��C���i�]�|	�<��Di�W��j��ZE�D콴����8
j�❳�x5Vٹc&u��3u���G5�%jܲ ��m|z����<3?��N����y��P��"�����I�8��$5�^�t��<F3Y�7^��Ae~^�����iJ�%���VV�kB̧�IP3'3Q��kHj~�MJ��_�~��#�q1�'϶&zE8cکc�x�_�����c�F��cJ`ʎ�-;�_�>~~��ի8��u���މc_-��B��[���O>�3��$��yG��WL�R��2:쌹�k��n.��%�_�d����kp�oB����=��������:�I�XA�� >�����_>�J]GA�1m���UQJ5q����/9�~�Q�+���{��w�};�v�W���?�8��E
G`��?Vq�ׯ��S�L�ę7�.�n5�s)��*}t)��>:���lxV�UB�,|g��gɽ�e�`r�B)���Bg�v<�s��!#�������p���"��I��{�ړ<=It!�w����������L�S�$�*U�$�.��\-��g)�P��_odz�'St �@9:f�ʂ�֐�u���W02����RZD����i"�N`b��O~��شD�&���᭸��;0�J���y�=�Be�3����n���\�jS���x/��I>l�����+���	��c�1�ҕ�����:�<���)���`��� �e�(�Ϡ�ם~�~��(����Ȭ�K��r0E�J��f�����G��?�G��xx��]�j�q ?����ԉ�ղLb�<G#�VQ�=+fM�b�5+��A7KiGD�Û�	aE[�i��2��E��{zɘN(0%c��T�.Z�W�����SsH�����w��5��'���5F�t�2]��b��}�݄�w�#�jttT�v�ڍݻw�]݅S�Z�O���wHS��Ha��Ƿ.�n��^��.JU�8R�g��<�/���O�WU+NtW� ���ߡVob�}���=55��.�?��嘝�B�^��2�\��D�A�T�L	�l�Ҩ�&"����"��Ɨ��*Š�F���T��t�����c��SO��X���44;=<��I��w�cǞ9�Il>h>y�;�i�2��u$�u����\�'�#_��RI{=m��=��7R5mSֆ�Ѝg�xd�h5���ج��e3gWig0V����`� BD�Yf<���Iu�,��n8n �yM��9��dEsM��k�j�U�[g3��P}�$)J�M�!G��&�U�"e�b#(g��{8Q��ާhep���jN� ��R�����^(�[��1L�,U�~���ç�:��8���͓�'ўWd^d����s���P��Z#]�䬛:^��U � �f`j���_g~�Z�� "�hL��3�������FP� ���)c꿼�^׳ߨ�5���c�s�TF�_+����F��O���!|��4��{�(y[�R#��+�3���F���&{��V�е�=�QЈ�_c`�d�{��jV������j0k`k��gW`�+R�;ϰ�{	C�-Z�t7�9�^z��H|���y9?|sn��#�[�6�!B�h�%sO�s�6�X��E���h��g�9�L��$�����zl8ۀ頰�֭W[:󫧋�*Q���{-c�,F�J1.d�b�qcN���^�����Na�[�<�K���¼�d#u���b>��,�L&�a.��e�����⛑Avl�\F�C�^�`TYX�W�G#��|#�,�"c���ܜ�';�R���atW]�B�ϛli��s�-��5����ʵr	i�����X�muK��9${L鸬�i��� �9��G�o^�\�yW�,�|��������ο��p�:��y=>�ѳ�1��_u;��`�֭8��M��W��W�D�+�ba��6���<��13����}���0�,�Pyt��u��"���o�+^r���Lɘ~�_.�7?�Ś��2^&���݀3��<�}�qMY�^�i�	�\��{z�F�'&p���@{��>p�ov��ހ��=���*��U.��Q/@�i��D=���4�x���3f~�8
?<� ��C��m��4:(dzȰov�8N8�`���	q2�U*x�����o��T�\i�B��!�@�*��3h23�`�V*d�v�jLL��=�[X��=Ә�]Ы��T*]ޣ��8���ÜN����%&��&��	�S,^?{��4�H�G��%PX I��i�Y�[a����>�l>x ֮]������o|�g�����ϢI��BQ��҅<rE5����4:h�Wѩ��d�@���;�V	�&�z���}&��j��̩�Y�V�12:�b��rJV�jM��Z\'fdef<NYu���ɶ�����׼p#�L��|ɥ͟�:ڤ��cjv{�f�}�Nl��$x�1<�s����0�
�u��_�V�rz8s&e��~�� ��TwϠ]k"_.��z92e�r	��Q�	�U&�����RL9.��X�{G�:S*#?>�~!ZE�=�@I��yϥ�OH�ksj^�iNz�t˚��J�>q1�qKp�>8�v�5X�b���7�]e),V��=���ns�2�����5@���tX���0�X�"�|7�vdR)�Q.�u~����Z�*n̴Xeq���������ѨW��vP)��ĵ�a�	�.K �ˋ4\�oSi�u����5��o�2\�ѳ�������#:�&���7�CTs?S��]l�q�����~��;��i�J�s֙�äJ�$_��K�����G�WBy|�1�~�l�5�����dF��0�q�[|��ux�������ͫ��K�=�qߕU�͡Y��1��S��z�2^-h��o�M�PDG	�s� �El�1����ɥ�6��j�$0����9"��KM�x�u��Q�����_j d�Ɩ--Mk=��}ӽ>��K��)9�3͞P�\P_+E`c��^�&豼S�-.]�Z�kT�eI�0��Pv[�e�z|��ʞD��6ѝ?%�;P��ٺR��I�]CT�	��� d<w�`�'b+Yh07z93#ɱBv��A��������)�����\��}{�O�.��C`!����a�?�Q)�	��-7�b�E@~������$��1��n��l�2W[������%Db@l�+�T�1t�Z4��|ϥ9�O��=Lb�[_��xKy�f�('�>{��r�V ����Q'�s���D} n����tmUW��${�=��v�u�R5������ٯ�Ak�b��kg�Ϲ�g}����$���|��g���Yߧˊ%g����9�s�}_lM�t��b��(Ι�JdH�k".0���ב)%-��"Y��{D�1ulq�~W�;��M�Zm$
y�	!QA'���t�������(q$a>4[��Q����f'Ƒ#c�T���jJk 'd�x1�ܹ�F�RC�=����t��r�<Q���R{ֽǔX���e8��U�xr���#���?��a\�Ky�|�����~-#�:|���>�U0���w�+_�ߺV�O���N="2R�*���ֱC(.U��&�8�Ԯ��a|�����N�Q%�j����LՑ���}+^vڱ`�fG��/\�_�J���~+Bܱ�$^�W��-�9�T��tQJ[��ж~{&�t��%@�6�ǅ���۶���!_�lKJؔ�ă\x�F�����#:��C��;5 �M/����q�e��L+($[�@�!.f�P�Ɍ8�&�4��"�Ψ#o��Рtk��V4��X>�c�y4<`_�U�0u�vO��;���'vh��{g���xcKUI�����6^�a�%������ǱFj����j���S�PܽXfEcU�<�Rc?�ĵ)�3�bQ&��KR?:��n��:�o�P����0�eehq2�A&G�<'���VOS�/R�#M)��3�9�𙖈�< �2��q�H�WS��sF�FQb�H'ѡ+/G�4���a4����^	�_(�x���%'o�=��A����ON��;�ǽ�=�m[�c��a�펍bI��O!�-���+�^����~a�dM�]��D,�d�+�iw���{�f�x��ªeb~�%0e�'��A�̽�1E���Ԝ Szd�i��G�C�4�1eP��S U�=��t����7,֨*`H�&.Ʊ|Q,���֯������6fgg�0�3,Gdl�|e��J�E������qְl܋��q�_`��i�s�*���K�SqBqvSYhc���0::��1�!�$����k�t]���Ѿ⒔�4}J6�ҙ�6��ѭxd�C8��ga||D ��t�L�5 �4��~�K<�eVL���3��M�K��)<���W��O�G6B`:>[gLE5�3�,��f�%�����R1w���h�e)&)�W}#7F-9�Plɢ$=����a�����b��k-��C��n,��$���kǪ�i+2�!b,�z?�� �T��Y������f�2�3�':DL�% �u������p�%�L�v���:��hsz��\s�⦛GE����0p�,����[���%>|�[���x1��Vɬpj��:{�,�h�E>.�R�7(H��Im�!9�����l/�yҴn�7;$`M���:��z��tˍ}�:�c*,~��)~bid̺=����E}a����\�qs�;,����'�Kl����!t��N�����qۊ�܊�ՈO���&��,&,�kr6.yR�E��\��N�D{F#�K�������`�wUy��] ��	1Q������}�}z��=�<'t���Ǵ]G1Y�s�Z'�t��QG:0�&�G���E�K�A6�l��~�u4�E7³���S��:�U�j�G���x[��[�EnE��)pA��2H��j,�&���n��i��)#5RF�lg��3� �CA���t��"�n�6���BE�K���(rc�觵=�YM�ϗc)S2�4�����n�.��>Sb� ��i�fEA-�j�ќK�W��p� ƴ�d��e�
���#��)0u�

���>��C;�����~zݯ�};戍��Gށgl^%�e����Wߍ�}�'���N�3��/O��z-֭(�"=��q��3�/7��}bY3�M�� �-�[�߸�߽�wM��P���DbEӏ�/;�4	 wT)�7����d��b�1>�����7��X,Q`�_�%�[��D�@��E��#�c���W��[߿ONw����8�SdW~��T����L�ܢ�/U�h��N�P�R=�5�C�Ԡ��U�5��(�� gT�%�i5��R����`*�Wi�3�~�$L~)w�,�L
��t ��&    IDAT�306ʱ"ma�:��L��_�>�%��XJ��\A�1��b�R��������'8�j~T�4I��,�i�b�Z^?W��FgsY�"(eჇ<��l�i]��� �^3�4��Q��X�o�N�L3
Ls%t�=���4�hÙmO80�k�5�<%0T�;D#��N�^_�����#%����qTL�ّ�d�H5�2)/]�9�4Ƀ��D�"*���i,/sFf�zS{���'�ض��.�E:/I�qbKe�I8�+ �/"=����(�لf�,Ba���e/À7��7���*���Zl����z�0��B
�$OM���J�:�y�%�I��g�JU�)`��v�G�R�*k/.'�*�;1��J[F�pl�����:0ձ&~���{��G�RV^)ٝ�]D���C� ��J�g����vƩ8��Pҫk<>�}5h0c)�1T;ؾ�qlX�+�(a�ޔ��O��j1W���4�-���$gbEq�M�n�
����A���z[-�����p��w��c�Ʋ��#�n^>�f:���w��ƊY�������ʲ&��ׁ=�J\~��Qk�D�KC9"a��������#�F4_6`�ʞ�����X�5GT )@ֿg,��E~�'��3g�(�>nC�����<�.�̤���wI�'�.K�����FW��"�d�.#s�-N��T�>?����Ig>Tf`ln<E����]*&����S���h��5�q��������T�L%��DF�������N��yu��OT8��5����,�s�ܲ��BY��'M�ԙߏ3�g�yb���GՂ�%�J.;TE���@UU�$���Ub����	��@�c U���-}�&�5`�%*���� ���q�(x,����="�]W4��	sg�--������8H�-���o�/a\��X�e�;��]N�h.��D)���Y>+�kĽ�{c��ｐ#�Mrs����ʁ�6���Fθr�i�N)�h�2DU8�9�m�#��\�|�� "�8���*�h�jͶ𜧯Ň���"=L���o>��=��W`�>��Ǒ},r���o����b~+�d:�7r�Z"n�h�Eԃ���`��%o^4dn@��R�(-@�a8��ը��qJt�%�DO�z�sҢDP(2ܼ"�ꉠ�'�D1c�C��)ou~�vG���(�##���'��+���u%g$0%��\��i�RL�+�i��T��^6���)�U#�4zf�Mj�c��
6N鷑��0�X��_r��ק`��E�|�k�F�����7LoC���чmħ>�vs�*��$.�����o^�ݻ�os��"�~��q�KO�X��z�yP�� ��Fm�-n���.JO�͸�Ƿb�A+��̔l���g)�E1[�?~�,���cu�@`�_�.~���htr"	�������g�W��x���A�w���[���V�Z�gs&X%�J�����/n������v�yq��ˠ�5tr՝[සU�Ob����YL�=Qi� ��sX-%�5� F�W�d���x$6���E��m<��#��0;]Eb�h��4��9C�����h��r8��g᠃�C�ݴ~��6=���o��ܹ;��iE�FUX�Ď�H��^\��W�R�w0�=I��Dq�h=Vє�Ȉ��y���?�d)8mЁ���~O��ǟp�?pLLL ���m3��/��COV�I�Ф3g�eR"���!6K9dQ䴭��������x�K��y�Mٞ��\�l������>r�"�&&02���>������Ȉ)}e���>� �W���X]���,r)�l%�j�eh{���F	�e��������R�bQ{#x��Ɲ[wc�Lu���H�1ƴ�`ڙY������h%�
hy|�vf�)�u����%0%`ͤ�b�'kWT)/M"c [h2�� �X��Agv�Uʖ��Tg���c�_\w�׬߰��&�XY�c�?�z��q����Ꞁ��Yn���9���?������nÈF��X�N��m㑭��������n��g��+�GU�*�S�s��ǎ'������J�@��ʦ%�b�  #��FE%�jZ�akP:�|�	0`fz?��Op�)����6k��Z>0��x����G��P�&��<�3*�M`�d��W���W�#�ttr�c�V~c��*PP%����"b�0	U'S�Q��b���+ �Q��cx��c��H}-x����x��0`�ω��/�9;2���H�i*��QSd��٠W�{��9uv%t�ϟ�K)%8��4�s��c���ޘ���0�w��|(i��2�+�g_���DYL�}U���!��X��I+
y"�12L���â��lZu������A\l�T@�Z�Q��Ub�\3HŢ�N�4�wjE��C�͎��p��{��$�R����Fy<���._6���R�f�z�a)(��*v��EO�=K0��^)�����Rp�P���?��[1�"��^x����AcI�g�\-�A^�e��~���)b\�Δ��ey�?g��jCЬ���&ZA]M��@�cy��/���?{QD���k����ǰ0�y)�MJ�Tvu�V����S�0�	4�6&��?h �V���ڭ*ʩ:^��M8��ƾ+S���'H�m����_�#W�����H��ʩ��d�/|N���4���}c�C��j�w�CJ�Q/�>�8�x�9�,`9�'�K�����5�y�	,�͉}C֬߀��_��V�avn�Ni���P�I�$������g	�Y��n���қ$;6"�C���i��d�!T��ǔ�4�1R�"R��l!K2OR�4zYcj��~��Vq��jW1�\ě^�t���S0J�O�c���)�߾�}���[��>���p�!+�1�M��?�����صk�D�l��
�}�_��g�<G��He^&)��������?��zb��@���'��^��
�7�Q*��1F�UC�1��`�l�;�l���O�jw�=�㗷oW^&4�^��p����22�*FJLm{"+��شi�}�Q��~�N���Q\z������^H��3�ĳ�I���B����UhA�N��A�<������Wy}<g���f��h��G'?� ���/����_l㇗^�+��]�����$ ��S��M��8�����E>O���@α���n��9�V��2��I�;����Xp���R�g8��a�8�hß�*��a��`u{�����&q��]��x�K_��O?ccY��-�s���q��c��E;�� �G���tg�ee=d29���8������΢��1�d���T���d"�2��TWlQ�ѓS�ԌONH�c���h�^k�Yk�,�T�@�*��1Ege,��={�d/|�8��Gaߕ9d�nz=��<\�}�t#��8>�,�|�z��*����"�k�ō���\���ל)=��r}�#��,�Ֆ2���#=VĠ�`*�֌>��@�5��Tk�#=�U����̮�Q�y�+/{/���Dr�֟����uњ�CFS�_z��G`�ꫩ�ҤShw�ҋ��>�os�]xr�n`�c��;#��?�^�t!�d��y2�5dQ7�}�N`���\6!=��N�Y%9n����v�܃[n��>t?^t�q��{ފ�cz Kmj��B�H����}��a=��#Q,灄:rh�*����k��)?_n ��x���n[F"�y�����o\�}��oz�[�g�_���5HJO��nz7��>��������Ƒ��D���Ͽ�����4�_���10@q��^��������(+L�͈�1����?�w
�
�B��O6�L��� ��K��.HJcpj�ܼzm�șХ��!�剼�Ԩd����x-4hr�rY?W���@��O�>X�0���F��)���LG���S��m�<�2�fB��,���7Wٰ��KL����j�|\�U�o0���cì0O��}'yvVl��h��z�yݲ�x���0$���>��W�׀�wu�7"V�eLV�PHbq���K<>��Dǯ1�A�S ��x���T���36�J��@Q�����₼��Clgx�Ĉ�}\\�+G
?$��-��g2�c� :����Y�CLHG��oc
�\��_��H�h�H�ڱ'*?'����Оi-������~	��sIa��n��c\�?��k]O�LN�i��~�%S/��ʗB���E��g}9{�g2��`�A��k P]��Ћ�9$�T���j
c�i�D�����Ǉ�y&�Y��#�/�'��w������ʻl��3��R`�
������kHn�+��@�scc�#����إ�~�"�'����}���΂>I�V��G�Z��&8p���'�ʤļp~n33s�F�!0�C�}�����C���P<�����@����yQb�y?7:��Ӟ���qO���o>WS���[�Ii�E�5��HI�i;�P��̝WO��2o4�3���tY��7���٠S?+�7�����i&�0m��8��M���a�t�9����>|���{O�)��Ҩ���8�o��7��q�J�6��Mp��Ba"��Ω�ʟ�^|=��J9ZNf�1�k�k��ہDbA���?�n��9GF���
�^��nߊ�ZB�ܝv��]X9����Lร�	��ukW��f&�U�\P6!D��t���;q�7�=��͕�͗��*b�q���͒*�'-v�,��Ƈ�J�l���i<a�:�7 �k#�h"7X�i�����/0��P�c	����W^��|�R�:���q!0�j��1��]\�j%�-��^���lٺ{��%�s�B:���o`��������4�j QF��Jh��IS�˘ǲK�{�Z ��'Z�	��iU�2��:�p�OBֺ�g���܌]s'*�<Zd��#���� cb�D� ��`�g��l��0�j����x�#f�����������؀3LYHc::>&k�{��j�!���v���VP�,x '���tZ�u1>�ś�x.^��M�̙��)����rIR���ZQK�9��Z*���7�����q,F�&0������&ij`���=���ZHSֲr�Jy�It�d۔�I���U)� �Z���9���Y�򖐟`1�&��=��>͔!0�Y���ueL%YO&mά7�h�;����[L�֬[���1<�c����l�j��sΊ� W,�PX^K�A��"z�E��Z�%�w���\�D_\�3�\���4*SO൧����L�)�b�l�����[oF���7`�ݸAY``/�ˤ���k�<o)Np$�r�4U'<)��t��c��_������\>�QM,��$f��O��?��. �o��b9C8˵E`���������F&��<>�>�ɔ SIl�HzkI쑅�6R09� ���^Gh^�d/s�`i<�H�����)��f�d�*�o�)��I}0�I�\Er;K&"-�ǈ1�Ri�3�[g�&����>U\8w`-�;v�
np�(�Z(*�X�ɍ 	����h]+�1�ז����I>�9����7)�3(�����E5~�Ck@'6�љ�"ud�iM��!]��E SUA�#:όB�B�ݬ���l�
y=�����;{��yDa ���C�	��S����?Q�����!��e���4�t����F��>.��k6����`�G��K�N�]���W����9�i�>.�6��x�j����:~:�(��+x+��y_�j��������=�x�
'A��c��K��%�1T��(cm8?�U�N+P�Q���D�f��m Ɣ?�`�n�:�N]�i��8?#�G�d/>�@|����>9��}���X@rd&�o@7�Q��C�֪bl���B���o^�q�>.���B��YwP/��J�+����3�}T�y�̯z�&�=��b�D�4�}8P�S���jU�L�`fV�)��dL��Ҧhq^�)u䮚D��Π����Ą�R�~�+R�\�,��-h})<1/�ď�\:򲏗���������9N 3VB��`J�4Hۦ��&糄8�9s��9�<;Hv�H�+X���-/=�|�I�30������R\��^{���}�>�c��V��p����#���03�6!�e%f�LG��:�y8���19J�a�\G'��%���>1�ܷ��|n��w�PZF���t�bd���ju
��Fru|����i�Ky+�g��]���G�P ��Ku�1�u�Jx�+��?�xl\?*�<@��x�F�Bs�����~������n![� �y$R���� s����0�?i�%��O|&����E+�"I�&J��g���c���F?��J��'W�׳!�L#�k.~Q��$�,H0��ީ���d쒜����~.�V{����Ac��5��-��сɏ�)��50���a���0A�;e���E6�7��L���KB�
�)�^��{1�N�|�~��;ea��yK�)�4>�ff�"�N�BJk�����P�P R)�9�	{�@��{ݮ �|����1y>\%�f[\y�զ Q��12��1�s�ghw[��d�zx�N�+NY�+Ȱ���|�ތ���}�бb�@[��?�?�k0�6g��I�Rs����"��5;�(��Dv��^������!��'k �&7h���ܢ0��nO�0��R�Y���L*x/�'�A��G��Fkj��*'���L�h�R^MN�1�Z��q��������">����̤�)�B} 2�m�z�)��X#5ڭ�2�r�{]_��.*S@}�|�1��;_��bX���NX��A�uˣ��7wb��e8�c12F)/כ2��fC����H?ՑX�py��Ğ�$c\�l^.)�x�G���/1���'>���˜>1�I�]9���k������ �{�Kp���H��6������p��o�b-�ʸ�����{f�52����fN#wǊ%XCFN���]=����ZE�ɂ�SŪ�0`�(���t)o�_3�q��LۿK�3G=�.��*��i�`��m��֌�1��ʞS(� zϡE��b�=�'ax��GE�Ȭ���%�ⒾD#����[E�� �
�!�е��|J4c�{����\��)���?���ʙf.��E�=��i*:��p��j�Tb���[�D��+P�&V�s_��#*�W���/���JA ,Cʹ�Lr��(DGn&RסN��m�x���/g����3�����k0`�tKJnE2j�*�
�(�{�����^[��*�{�_�����͖�~N�`��ϓ��?C#9Ql���_n�&�{<7��%J�pm+�ҿ	�(����Z/���rӨxc-��<?Ⅸ\ޞ�,5�Z����7�B�C�y-�{���ST�ek\�x��)e�\�t��T�u�5�LO:z���ϲ�0��L2��g�����y�G�bl�:���H����G7�ۋ�K�l_[��v�[�7K[�H���ptOD
�Uj��?��:�fL{�a4�N*�G��~!D�S�V0=;#R^���f�ǐ(��M't���4F�Zө�Ό����Cs���BE&7�p�K��=�dL��ҧ���#c�*�%c�3`�ݝ+G�����^�� �Qگtm1v�'߾�E�ې���ӓ�g`�q1-$�m8����U��*6��<b���;�Vȼ��v�^�|�⛱sw�x�S��*H��Hu�aE	�=�h<�cq�kQ��,p���
e���cW���\��;�}��n��z7�\a������YE����� �����S6GRޝ�1=ﻸ����_Tƪݮ�T N<���3p���J%u��_&��/UK q�4y�E��?��]};�+�RE�"%��yP�%AhX��J|��&��{4�2-��Ɗ0��A%�t��"�r�&&
|�Co���K�cn���s1n���z*��b�43:$��X���E�=E�+�{jؕU�d�6]��o%r�
��KF9��R��W�KxJ���������J��j�+��V� {��u    IDAT�>CI�T�̝P�Y��1(���z�	x��/ƚU�vS������&���?a��B��;G)o�<�@�T���f�!�@�>��o�>��e4����Q�c<��1���@i���
L�~��&����28�x�6e!��6��~�c�h�}�K�W'/G�k^z9-����}W������5�zG&�'�G	L��=��g%���Ŕ�C���4��tf�z[����eR��h'��M('�K: �v��Dn�Ū�&pflv���hY��ma\��H��1	�'HwHT[hO�#I�:Z��u|��$��H��^�cB����&�/��b�*���N����g36���>T�piR�j��D�~�lf:�
t�h,�A�3��<�P|�3�����	��hQn���}��X�v;�PL,�[YBm��]��B��R|��f�1�hW/�:�ɖ��%N�>����\���E���Oa������ȹi,P�q�}�ٍw!��]o�K�yK�M��������4FɘN,� SMy�4��01�bO$�du�%�� :��q�Ѿ;5G
`�cA�iI�0Rf��`0��^��=���x�zL�o�aR��ؑSc\���[��JeE�B[������JQQ���d�a ��&�v�V�үu�%>��q�X�K�WI���s�=�
�C�J�j�iq�&�	ܫ2�����B�K��p��B]��%�C�eO�n#���Rh	��%�&��O�%!g�`��Vf�"�D��kߋ
+$|+;?eN���3��E�U�^��f:)��w5n��x��\&���z�$��ӕ��ٶ�S�{���HfH���;A�&ς�|�a`�1,~h��o��S��'���YXaK�����v>�s�b��|�,)|�k�b+�nܶD�6��Q�L��N���i��w X#�!�X0�.������y�U�@�ܢ�0���t �oz�`�@�ob7i�--���hĎ=���9W�"�������{9�ۜd���Uo�#K�)���)��=�nc�*l$/dq�E`:����w?8���:��Z�~&+R�v/���M��"Lԗ-�N4G�E���qEP��=��Ay��/5�g�4�Yj�TF��C.��3u��G1;��D`r|�n܄��q!+�8��J�VG�3�H�1�$%���~S�7K�yC`J��Hy�%d�%$r��1����{�%�5ƴS���RƔc�Zf�c7���9�&\����- �U�����蝯:tI�o{L[�ހ!�1ӯ\��~�l��7oĹ�PʻR��&��+���\|� ӑ��ȣׯ�׮��Z@���T���B
kWL`�M�z�J���I��j�V��O���=��[h`�ʤ4+,i?�� �ӊ}�N�)u�Jr��BL�5��g��N:$������{��o�av�&.4Jic��q���g��ӏD�Θ�‒׾8�N-4�kzV�r)��+�QΫI	s�Gv�n��I�edEID��K�V��1�
���̩01�9�U���dA��f�d$h�B�B�H�inf6��T���Y��:�nX��Rw�q���q�t�4�Ĕ����P�]m�\�+	�:�^e�IIX�Aк��&i/���ɨ �R��,���&.Q{ETf��w��M֒*av�0PY���V�59�CM7�ܚ���+�jR�4�+� ��6�}�M.��M`Ӧ}q��c���9�å�_�{z�>m�H���EJL�����E�VۜQ)U��Y��df�K������%�~M<�X��Z�ϋτ�K)���К����i��2.&-=������~)��Epښǲ�>�z�_��ǭ���'v�1!��:ՒT�-�$����l�L���ӻ��PO����"C�3�q�����$Z��h�-�L��5�+V 3Z�@\y{h��H�&��SY�AJQ�M��ѡ�y��
0��Qb �u
JY{�q3�V�P�\m�5��D�����ѥϓ��Lm�JS�f�^�䪓�A�(��ȳ�ttȴ�wٔ�� �%���0a�S��zc�'��O��"9t�hV�����c���~��������ضe~w�X�l�y(�'ǌ�v��.��:����i9��4�����j~@�I$�y��o��5|�����w	�gg�O}��4L9az�\A`z�]�c��7�O߼R yk���+0͈��H�l��U�46��Z�/\��7�4.b�cXbp�Y��]EL�%�^r'bh=���XR-)%���U��4c�dȹ2������*��I��߲�A�D;�2��a@��(��Y�j�̒�����ӟ���>�T�d JOr<�}�!�'�r���H��+�&����K}���a�1�_
VxlvP��j�t�f����=d=dP�x!��,{�Z�^l��N#�� ��K
WRx鉪�a��-��஥��ԸL{���2Ę9HSō���x؇��M�*�tL�R�:�)��brDd��N
?6�Z7/%~o�K����0W�p�.=��?c�oW]e����ky/��D� HU���T{E����Q�QqDAE�P,�A@D@�� E��Bz^���[����9�>�����	y���=߲��k����rrֽ�����}�R]m[�F�G�P<W!q��`�W��t�b���qgi�T˓E�`BPj���v)a�N�>���+Lt��U~�Ԝ��v��C�R�R���̏�& ##"-�X��@�s(TӮ�3ZW�S�F%�3E֭�_J�$Ya��q�w�`��xY�{榷�ݘA9U�ѯ^�ϝr� ӌ<��X<?���o��'g��#��C���I�Ĉ��[I.z������g���ֽ$���&Q1H�&-���Rb�*��L��"S�
ev��
H弬��
0���Xy�-^�a�m�V��/z��B�̼�1$Jyt2l!H�V<%yjp��YI坮H�I�y�th�lʘI�W�PVE�:^u��::�e�R1�`�(���ᦩj�L�ZP�$,FT���:�1=�m���`���.�T^f B`��ۄڱ��;(0ݍ�G�d����p�ŷ���=����gA�&��M��u�
R-Њ�<|Nj�
;���ϔ�ʖ�Jt�U���F���
� ��j��Z1��p����^���uiRS�������g�qK�f�D+wY���˻���w@��K���]`�����+��#�LN"�M���^���P��J�X��M��'����l(]h\��Q:��蠴���j�[	���1$�R�xjV*nG���$���Kv�mN#��x�02�6nX�^�D6�,u U`�E���;��=Ӯ%xL̄�2?�2^�j���-Ѥ�\(sN�L��F��(��M*v�y��1z���M�:i��%1�7Z�1�k��ܜ"�k5{�B}Vԛ���;=��"�D��FGǰh�����X��&�+mV��J���bM��L��B��J�Th]ҟT��ܬ5`�20J�L��ƍ:��Y)2�ۊ<�>r���eO&Ѩ���ݠH]�[�t�B������p%S����u	^��B,*�1Z̡׬!��jTP,e���{c�D!dp�ݼ��'�|s�R�R�<�C��LW�� ����c��C(��q��<�u���;��6ً��t��hL[L0a��^�H��1d#�ZS����h&����w�L3$�H�PѳiPn^��J�9�����c3�0��a��9������@U6`ʩ
��ŭY�bz�����L 0�D���u�ZM��[�&�2�$}ͺ-�k�H57��\��>q��W٪'a�l�,wie���V=�r��}��c�l���HG� S�'o����DF��L	�4K ���R��E5�>� ���
Tku|���`����[�����=��y���s�ˇ�*��k�����ߌ_���TR(/�������lF-W�gc��(�*l�8�&�){Ņ�*U���\F�<Q��$C�[�2���V	��eu�)��ٟ�].�0�5 u��'C<�����m�d� �X��.�j�4�v�	����?"w��<��?����e􁵚n��sB��l�������CT⯳g�T�(^S,{̟X�r���Zi�b;�\��E�n"٭࠽���'��3����>�k��
O��F��C/���S����d��Fzn�#�I_DZ�J�u1I'�u͛�dy@-A���&iv��U�Qas(��ը��n�ߩ"�jb���C�����6W��^�.�v��1��y	p�$��<rΊ3��%w�o,!b��'���I�a�iM>GI���	���i����z5x+�(U��^�/�1G���}�
7ms�&cFI}��5h��Fy��M�q*{E���&�s���G�G�o�ۮ����f�`�̱˫�z�.�iy�Y!����%>���d�ǅ���2��*j���1
�=��|"M�,�.�f��/�p��c��?�xl7�@�q� �i��S��=>���2�/E?���0+�n:%k����(S)
I*V�6��z\�'�#���$C�H�E��:��:�b	J s�=YmJzZ+f),(��g۹T�ZS��P�5"��	0�ƴ�"0��\4ᶇ2O`Y&���W��\5��R�0e�%���Φ|:%U�^��v�&��K�^֑!��t�	1��u����q`��%�+���+�ǎ=����X��TH4i�o	�kg�o�s���v9P��c�������k�//ъ)�4�d{ ����m��/�R�֕��Y
����9#3VEY��	T��-_V)�&�朥Ɣ�[�2-�4hm6`z*^��A*�wι7��8�lm
E ٫c�����}8��@��	:���U7ލ�>�\lٴY�����7�+_��K�`]��/o����h�A�r��/�Y�$	�il�0��L��Ҹn!�)0��_�`��C��$�O�V�.{��$��N2<l��i �Zx������Q�q4 #�2D�!?�����d�ͅ�<m��A�T,����ī���
�6_W	�nn�qQD��#�F���FH�S���0�8��vp�.2ԨZc`~@�n	ՠ�H��M��Ϡ�E2?�n?�N/�lvH�(�.�	����u�N2�$�q�/fD4%��t2���S}���u���$�����W,�&0�4VՊE��lY\T��]�v�V���@�P����R�E���\�贅t��<�����֯E�1�Fu��y|�3'�ط�����I����7�_]��J���짺���-\�-�f�it2l���5,�T\�	w��ǔS���ȍ��bJ`*�Ga�c4`RN�6LW$�'�8j9IMq`*Z%ڱd+K�������i S�De�,i(�������7y�z�+�E6_	�ئ&��P,	P�>^�DA
��B�s��ju�F��c�FOR0���r��^��V��o>dW|��ǣl�4�̰,�[��~A�9<p�C����eX0>�5�a��NM2yU��Q�T�xvK?eV$���g�{�g]u/���*,�qG��}���ذ�z��1�W\� ���(dR��G��޻-��,�����/����혭�Q$&,��RO�@ELd�Yv�_�U�"x�E��И��@�&��U�=�N�h��Rא�՘.��FӫL
i֎A� �`�a��iu�niH��56�:�4������PX}r3�AM� ��ýZ���g=�_5�@�(*ѧY�����F5��|����6���xp퉼М�>;���uAx.["ԊkQ���V����6k�j��k�I��>��#�޷�!󭨴���������-�<����n���:jOً�됲�,�K4O����P�r�z�����_��44��4hH�Ǯ�45��y�ݠ�n��nkC�6�<t%>��7c��l	-��F�Sp���8�G���E*U�(-��o����q�p9}�V��l�=�y)(�錗J�x�ɶh^�Z���&�%5���8t@�#O���~��$��N�7�e��P��&��D:a ]A|�X%�"@5҄F���is�uĖ��I�����m�(�ǒ��~�%�O.�=�t��RX��Ŵ��A> �L��y���R�V�c��=#Vt�����,�VfЪO	0=�������ö�Z1�V"!��#������Bal����"F��M5��8VL�"�=�^�^=���s���v&�u��{(�2�O�lT1���D�hB�G%�H�L��I�ɴ�,��O#�U4�n4Q��t��z��d.��� �N6):Z-JF�va�QcJ���+/�i�C�_
���̩���)w��1&��s��s�i 0�B��E+�WW^7Q��D��%s��W�+1�t	�ȴkR1�?SjL�H��9���W�x��$�o��Z1�ƴL��A{���6��\G�<,ζ����2��[��j5��)!8+D��&RM�������57F�r�6������M	���t8W7*��"�i8����Ϸ<!:K�߭ⰃV�_?�~�rX�t���[�=]}���J?�^������m��Hx�����p������G@��kZ���ߒ�30���`FW�l����2[!NWb��g�)k�=��&L;ȥ;�$�TI8������f�z�>�CW�]��=P3�N}�V4z$��Q~hL���U���;?[7M�g(PK���1�HC`j�nI�ĭ�c�	��I0о���5������c�6� I�I��B���%�2���L]���fE�ĬW>/$r����F�i6�E��Wzm�!4V�x��L�vn��S�~Op�X���i/�e��x�T75~�����Lu��G��2����D:����16f�'1�n#ڳ�hMmAcr#P��

%���x��`lX���T_��O��nD���e$�%d���ӎ�a9��"ڤ̰�E�2��S�VWz��f椱4����E�V誫�㞰e�.q�'=���Uty�t��f�.�fŵ�E�D���G
/��v:B�M��zS�?eR�$��{�lK��&Z�[��{�����kfnP���m2ش������YNZ�V24"��g�k����٩�@}�?r/���w������8	FQ�]<�����հl�2,Y<!=���K) uc��tf�'�-����A�D�C�Ze+�F �t�]�p�1�`��]�}Bw��82Ov���x/����8��t�E2�-2o:��q+.��6��3��bxlAL�_{s�*�d�%������{��5>��k�!���	[;���ų1�V̵�bH޶e�(XEK��[���Ӄ�~f�_�
��^�b�a� L�)�U�8-2���ˍ��8�G��<5`jUf��A���Q�m�k �=a�k����ZNr`e�)j�������i��kΙn|�k�?䚌k�P4ҷ{�/����[[�%����V,�����r�.
Li&� �	X�����?�[*	$���&2��A�ʁȺ��a��ȏ�|rJ�i�����N܀�U�9/���f6H�A�
��ucsH��X4��;�9���A�~��n��!�^� �]�ާ�����S�<2�!�X���9ޅ ��(�L����ϯ�E31>+�屄ϋ�苫y�Eyn�e�۫���!��q�_o���e
�L���ͫ��T��.3�WD#��Bv�Nu���kw��3y�sČ�AyD�gV��<���?������k�>v�=�[?)>3���'Qbی�_n���ԡV���t/suU`:�vsc��?|O|��o��a���� ӏ��Y�1-.������F&\G�Z-h\�q�ܫ3�����Jxt -�i�Z�g�����Z���Wdz���N�Z1�f�#���2L��t)�8��F�RG���u���Q$�Et�)���R��e�S��ZŴ�EujV=�hf��bA�ٴ�I|0U��߁)+����]��80%�M��1v��m-�7`��Z�hŴU`����G�?�����T�.��G�k�7�����N1��e����1�˄ ӭ-��b�qK��Je2��0 �����`�G�1&�G��s�,/KkƊ�TZ,s	L+s�mm�H��|�T��Е��2�b��3��TL�=tD������i��v]Vao"nB    IDAT��`v��^7���<��j,Y4�w��Vv�+�wRI<3�u���ΧQ��U+�l&�<�̘�Z*��tKi3��6N�����tj�c��U{��D�	W��=�]�ﵕ�K�i��y����6�I�L��uڵA0b:�i�����׫�r]�.�'��>���!�����M���� ��0ӿ��LX�Iې�f4̴U�"�K�2m�^)l���.Q�u�5��s�Ւ����|�:�pxЁ��k��ᗿ�O��.+�@�T�)@W��\6'=;��0R�u�o�+�2=�KW�[`��5�ìY�M)MJO�Cg�>��%����'h��ƀi����L�X�=VL�)�N�"]�`vv[�oDu�f�xLm��@0�R��S>xN;�CX0���ik_��y��[����ϔ����X��vK1����s��f&%b^���>�AW��Z3��M� ��ǥi/�@;a�T(ۑ>�YD��w�� ��ćiƔTK�ץ���{ժ�X0H^Ĭ��lyNT[L3�ΰ��Q�� )Mm+��V��&�� W&!�#`�͞�/���籖Q���ʃ�2
���\д*!.��f�Lm@��'�n/|�K�FQ(/޻R[�ă�H�Ria��͢=Q]^�
��m@ .@ѿ_�!Z�l��~O�,\��v�ʜ���aI�x5�O�[O<����č�N��w�@?H&����{q���H)�O~��cń��6��~}���_Pa�[(�<2&Yd12�i_L=��a���Z@��H������8
&-�Y�,�)��2�qmU|�:`�&���Hǒ{1-u��x ��N��؞牽xE#���4�;�s ����G�����Y,T�X�3F�u�Yj]��<.�D�G�a�?@��+�����J��	kUD����v樃B��u�B}�?��B	4C!u�D�Ԟ��N����'���X�\��L��̱�g���s�^x]=�JHd�Hf�B�c�KǗA�VX\/��g�m�g�&���`N�|��|���ړy�ЬWЬΠלF)Y���8�58`�E(�\e�M�I� ���Y�u��@a	���H�x�ȸ��+_�>�cX0�h��
�i�h<90g��80���'��9��V6Q�C��"�����q��N�1��łs�����o=����K�IF�Ɂ�Ԥ������!�ٍ�,��6q�u{;���;����Dk�h�_�p�ך�q�zM:z����Gy������̈́���v���m��N��m`Q�����~�����T^~�)���Y��)�'vBadBZ�1(n�۶�h�)c.a��X���ΐpl-����8��ic��}��#����<�LY�0-�ё�J���O:���(���0�Th��$��Ag2�`�*ӓ#���VXFO��}*Jl�B�%0�Vq,���.�����˃���%����I� 0������8=\F7�A;t���b5ug"U1�5�NL�.�SRy?q��8���%�q��? ��1}�|����n�K��Z1�(^��P;Ls������cӖ���<�6O�MU�W�����򫧛�o��ѝmi{�.�����wP��`nf��+���o����M*�B���-��1L�һ�T�ሃw�?�A��6�-l�b�Kӕ6�f�0<T��[qhF�š������≵u��Y��ji�'�v	4"&�������G��ݬ����V;���.�>0�ER��dR':M�]d�ڑ^PE2�A:#�Q6��M�&�~�=��d�xiud닝��EM.P��C�� pK�#�f{Io���-V75�Q��P&m�ib��,'�Ur�ܩU�� 2)�]���TZ\<�W��k�e�z�jvnV���N���>��\)�t�/��On�u7���u�G�"I*V*)F;��g��U�i�]��֫UM"0%mK�Q�J��k��	�Ԓ<z�+Ɇ�.V3y:�Qۘ�Jot�Hyc!n���eJ�e���:G��ii�Ԧ�۴�v{�z��U��5�S���ⳟx/�Z3�9����S\v�hݙ ��������eW`h+�F��������l#����,�FS�;C�"7JzHB\��<�u��i�r�j�Lm��f�͞E�Z� H�@]y2�+�����oiw����,�͎hW�f,TޤЭ�/�5�bؐҠԳ���+�]M������l���fO��d���w1MY>f+	�:-Lmy����������I(��T[���� ��m/����[?�g׬�ŢE�)2�"�	�f��G������"�Je��Z��j��f���cX�r7�,�g��ds3ULn�Ķ�m�\��ho�J��#W\wn��,+�'-=�	Lyli���N��7�Ҥ�u���2�aࢣV8L~�����5�Ti�MlFʕ��?|�	�F,��4�r�5Fm�#�feF�&� H��d����J�2ƣo�v]����V��,h4�6���'�<B�q�i~��i�����g���R���+��^��I��E#�I��J�ߛ꼢�O���D�ګ󁩞=N�����A(ea�ؚ��ZP��C�\3`�}(��.�A��,ƲM���W�}��q<��(À�!R�j �y��K������o�A27,�S:���놮�rDF#�c��4"dDUs��LS�%S�P���B��О��EEu��x�ێ�.;�Q�H_S<��Ίi���&~r������Ɛ��u'�1�⬱8�bc�n���V�*��TbBc	8X��2G��ס���{��-���כP+��ٟA�ݠ��^|o�
��Eo)CB��V��O��b��,�x'~��l=����`������2��3d//-F�v���.��L���}��[e,dDә����cVPuަ�d;fg�"��`�Ho9hg|�}���M��!�t�ԗ~�{ފ���CW*���ЖT��WF�*jT��=FL�WEm�d b�ƈ���j��y���~d�Dmi�X@"��X�T\�{��6OH��rd��>5��U�LiX�� 7<"��S��v��g�3O`�b_�AczV�/cK�Q,!]b�6-1�8��\BL:�r�-c����2�Fj�rh�:]ڲh��,�7<8��+�Ԙ�?�i�̏�j{�Y�ĵ7�-T����I��/_1.�E���檇�n�����0F�Fd0A��;)ڃ��+<D��r0��o��(���e#�p�n'T�I�N�C�=��B?<��8��]4��0=�"���c�T�DF3x����� Vl��V1�Nk�[�;� � �<�Pp�#|��_`��E���Mބ�FK+���U�m�7�@�iُ��C��e����n,���$�֔�v�~�l�D����עۭ���l.$P��C�� ���Q�� DzKi�S�\�f�Ɨ�Q$,������rpl�gqu�x�0�J�yD�lc#�7k/�A�V���͢iXu׌6f�n��$�z�u�M���Mt`%g���:�g���2!��v)~x�w���r�<���U��/o@?3�D��:�Y/A�ڷ��F3���Ԙ�����84��PYʭb�����a�#�CixH���v�FC��L-2�Đ;�J�c؈����\Iu0\J!۩"��*��nm9��������ő����r���;pٕ7b��)�o�`���0�1t���A3EWm��3A��+����FC��e�e���
ֲpv0r>1D`u�T��\M*�L�%�)����)�{)uy>0MuzH��Ү�2+�0 #H
N�1.��yO�=��"�f�b���8:֫.�GhYn�c[_/?����T�Y�O�-l��<�3kp��_���cɺ��J�b�FBJ����
�[[��7ݎ��o���K�.���Qd���ި�����MQ��@�:�z2��u�8���p�[߂l:����b&x��52�w�i��{���j�~ؤX��ʛq�]`��	|�o��;�K�R�&�KV�οs�<��C�R=��2͊2h�i�O�+�R1�LTBgIK�y�߉�2��D�Vu����t(}� W�Ox��>�JrXY�y�`m0���R�������+���<��(�������t�`@�%G��1�Wa�=x��4��SM��}��ۀ_ڼ�+�M��\�������S�4<U#ݚ����}]�3nG����V��댉M"��# ZU$�SX�8��{8Nx��(Q�:�*��yr6���ࡧ'q�շ��;�l���#�A��G�9d��a�)^5ƓD��$Ǩ�.���lk��v�S�F�">�dG���Q�c�����0At4�����$!:��i��݀U��G;5�F'#n��۔���1��gT�����������l̋�h.���~ڼ�M�Gܣ��`�/�&�^4�R�
��bu2��U&�@43��5��x��ױ'������{L����h��d��M�����l~ĿǜBt�c��yC�S~�졞5���w;����3��S�W�������^����V�A&��ґ$�t�r|�]�����|@�*Hb���o]��ܿËV �-�ɘj'�E�n)v��dn�Gl�y��|枯�!M�W�|6��i�h���	#S!�E'�BS�Ȩq�M8�t�Ow�(�[�-s5�k���ɠ0:&��ӖȕԗГj^�F��v������`2�E�RIZ����YŔ#��!���<�c�Tt�L���S�7K��{��R�0+9&��0*�WL�O��iӍ���K\�gRy��
���?��w\�V��.�=��m�<��pyD2����N�A�P�n�+�T�ԥ�L��V�:[#�
�4XF��� �Q���ֵ@G��9���<x�,���� �8�B����Q�'�/�P,&�r�B���7`��16�A���,�%�ݤy����ҟ��Ի�˽������MM���@��-cfV��Ej&=�w**�8�6�u����EV������������;Ai�~#��s�e��k�@��v��L6+�H3��$��i94�!�*
(�J��v5�D�i� ��B��ʜ�.������X�s��SD�xh���L��k��7fuM{�^X�N�Z"(��7�҈Udm�+)j(�R�Q��o�Q�ը�ܻ����&m�������f+��G�/|�SX2���V����}��ϯC'� �$Ai�jLi�$��SRy�Lk�o�+�HL���VE��2^kb�!�[)Qa4�D�^����
����상$�l�
�IYփ��D��7���W���%�H�	]�2@��¢E�(Ҟ͒Hl2WffaOP_�5�j��3}��'p�c�1��J֒�qR��G*�V�`R5��L��Nh�4�D�P`*��(S�XܣyУ��LU���yH";��G���r��|���x�i&H���ڔ�i��B�*I[Ͳg�����R��^�!3�ܘ�T�H鑖+Q<��gU������B2�*�`*T�d�v�[^@s�9���}p��`$c�b9�xz�Z<���XΆ���!����r�]��?���_�}���r������-�Ϻ�P�U�]��]���T(����{��vl�x1�� 33�xn����{12\Ɗ]�c�}���Ą�����i~��Z��/.�}�	,�v�>�x�b�d������.�	3�2�
%&]rZ��~�.�е9'��4y4Z���~3b�W3���t�u`�Sy��^oAaѪ� yx�&0J�5:��(�@1jg�/��%�Ile�XD�z	c��x�}����!��5a��(L� U�H����b�H�9�ʷm3���⏮(�����k���_�N�V'ip��������I���Eҙx���R-I
wh�8�nsF�M��{��;�r���k���F���dgm� �?<�K����{S3u4)��k7ѱ��(��f�/�>c��Ӓ"[ut{�c"��k#���p�3�u����X:.LG�P��A�T}�� �?���~�zd#*���1 �7�ÙH���U #0������g\�fN�P��N��,������FI��Y��1z�������u:E��b|B������_Ǿ�((������-�?�?S֎w>���"`=o'kX)gy�#�|J�K�/^�SZ:� �X՘j!�w`j�P@�$7t�KRT4�c�/&�A��D��%�I����p��_��F4AK@�sd�V���-n{`��;=������d=�CQ�\���>޳i��c�פ�����	��.��Q�u6J��1ҵ�ԋL�:0�AK$e*="���E���(��ijY��]��!L�L���	Q�Q`�v1h��bڬR���&�Ed�Jt}v����*�n�� x-� ����ʜL�̕7� �@�
����KČ�5�3�E]�jL?q�A8��CP�Ǉ6���_��Ѷ��:��/DcJ�q��W�w��cR���⯮x ����򎎌ax���;�^I�(-CkY5Qm?��6	�b����*�V�X
&H�l��ze3��$FM�����v�ㆿn�ڷ���w?�f'�L>���b��D>��P>�|�}�L�##Z0��Q��Ȣ����b�-X�a6L�Q��--D"U@���8�?� jT���c�S�uq�2Ү���h�:��+cU��Z���ݎ� j��E!�@�9���dcCYјq�x�Ҳy�V�y/�ۈZ��ё!���bv�"-<���W7	n��&8!aM-iv�P��a�.�)�Cg�ۦ�0T�adh�|�}��`��,2SM1hI���h�Rh���Uێ�;����L�U�L�x�.���b�]��ytH�$m3���^����f+5�[�&�#���~ w�1���9��x�[ވ�v^��T��/.�?��z�1d�Ȗ�H�YQ׾T�l��C�Qo�Q�!�1gZ���&�v���ra�gA�f�dߡ�c.�,+���� �.�{J�TTոJ��ߗ�5i�x�I�m�b�H_��Ix�@����ѺY��3�-���78����=�W7<�Kn{
S]>/לhLI�Iq���R1�5���.�(��ym��Z[��lR1�{{m�O~AȐ\cJ`�p;xp0E�%�4Yo
0%�X���p�qD�nI�g?-nÀx�u�4$������}遨m,4*/�5l�03�A���=���:�iC�j��K�������O�β�Q�V��-3ؼq�f+:~hS�%�P,KO�F��L�$}f�J�̑��9I"�&�4�B)�E��Mꖍ�q���Md�	L,���m����n��&04:�^*��7M��U�`nn;m?�����k�B�暡v�����9�݀J��l��|�,�c���Ae�+�1 �J%p�Y땭�P0��-^]�x�h�_אj�T.��j<e�J����J	3��Fa��������n��W�ueL���W��g�*������C�09e��R�X��!hTو`��K!�Αzk����ji\��C�KB�=��!1wIq}�lq|��ذ�H\s-g�]��x{��"�ɇh�u�����V��l����2I�5�I4g�aa���{Nz��pH��x�����O�*���+���?���&19YC��b�Y��<0��l�s����K�I&_�U/��p�0v�e�����ͯ��� 皨C�#_A�̈́�w��n��_������a�2�H��H��zl��f:v�*Ky)h'#�l��q�?f�zT�|C4��[r!����8bu'���>���5/�n�>��U�e��?9��rP�5�-R��yqz��ݼ���4��񤙼�ؓY:&�_�gu͌鹿��s�D���}N��=�p������a'{/��|����l2��V���k���Xx�.q���n�-�h1A��Z������ǣ�'14�:��esHfRb�t�� �i�4-�[�Jm�n���:���p��p����S�yH[��L
}j<�Q"�R�Ib���~_(��BОeų.I'�������9�E��SC����t2��*2Ղ�S3L%�ϳ�}T�1�eȡ�8���?��"��F��i��$AH�+��"���C;nD�R/�S���    IDAT�HѰLS͊�������4��~�O�����](������˧*0�>I������%Wܩ�ttJ�!m-�.�l)mkg��=ЬѬi��,g��z���e`VЬb��4M�eu��/��ڌ�6��Ηp�A� ӯ�Bܱ�Y}1�nUtZ�Huk@�!#�S��,�C�ڽbQhd�F�N�6&s(�.F'QByt��A�Ά��@$rpS 9O#(OL]��~,;ᮻq*�g�}3�� �k���!����2�f�C��g?������mX�$��<�"`�4y,�:�hS������j�=�`�8V�����j�$65,��Q�y5v�i9*�:�xjy�)Ԛ��~�쉥�'$�۴y��Ql�4%����7��9�UD���O��އ�h�����>po�|�
�8>���x�혥Eu�F>��[��Z�߾���������[-YaΉ���x�?���13]���ޏG�X-Ib��e��ð�>{���E��Ss-$�9�g3	��8��}�ӎK���KQd�� gl�����q�E���G2_B~hD*�"Zge'�#�o���Q����m�bm�<o���D��?2�B���1"}�ns�b3����)d2J����衒��#4��4�iMc�����S��2 /V�[���5J��v=�B�( ��z"����?���|���4��$�F�K�wq֝��E�F]�?��J�4�B�>���(μf�H�eQ2x-�h�1cT�N.-4Vj5��
牰H%*o����S1{���L,$¶��/מW�I�O)8��=�E����KL7.�ůz�80�gT���`:=���z��=p��NB�&�v�Z��u��'V��$�!@�M&�$b3��h�3��0]m�&�e��D�(I�b�(��J��}�%�M�r	�'�h��ЬNa|8�5ǩ��	�(��n��/��+���w�RB.���v�'��X츭RyI�'0��ҿ����\S�<�s�����F}l��C��>d9j��ԎI���k�q��i�B͚%d}zK*��k��cZ1����^U<��#�h���ΐ���������O��Jl��������Ӥπi\���H�C�*�;������_��C���= �'iy��l�����L�;J:D5f�����p|��}�`\�ޭ�f�t ���Cֲ������2s��k=j³���,V1@��h�ۤ~s�������W��xF�8�iU��4��D��XF��]����z��z�<�s35-:�[�̂b�Wbuɒ'�ʹ|&F�����_�W�7��c,� ��ؒ� ��٦�<`����$~u��X��T:|S	�$[F�#�
���"y�����O-{r1�S{���xe4|���a�7n�~O���pp�D E�S<S]j��q���U9���PD�'�*v36�PS[sz�ƺ��{L�@�6!����k$�=o�P���l���T� ѬR��}W�)��D¦���Fƥ>G��J�<��1���ܷ�ǳM�4z3}4�����N�Tێ0Q�`�����G�݈5f��x^����dK���<�sTn��;�k;lfs����Vk��v�����0���}��E)�}�Y2���gv��.�g�P�?IR���5zj�!h6��"�bQ�%jL�S��� ��؇��T�����se�1�b{��!�"�����<�%0eB��Fur
�&��ڣ��<ZI�Y�䭟�a�K�a��Ȅv=���pN>���1m����c3��w/�U7�&���}vſ}��A`��ו�u�waæ����аLڷP�i��L�1&Ͱ+��B��T�V�2?���jh}��H�*�곘�zhm�x)���s}�
T�f�ӿs�g5���,�v��V��F}�d�2ʧ1:TD!�C����쩪��M�V�X�v6N�04�١%HF��@W8|S�T6���kQ�{����������0��b�o~�Q��@��pN<V����xٮc�臎�n˲`�Ji�������}\��X��r��r1^���U��9?��I�fz����w�cE��g��+���M[�b�������2�w���
.����[��g�e��K�~{�L���4~����s�^y�����m�[ `y��9������S�Q��a��w�׿�%,Z<"�o��?�|4�m�q��oƇ?p<)�rm��>���v�G�]Û�t$>���Q.%15��~|>n��!��J�ͦ�x׉��w��w�X�sI�����M��wwمHf�(�h?�\V �d��
B*�u�=�h�������T+r���ւa�#�ĕڨmi�=A��FS+�r�R�ɈKt6�mM"n]f"��W.�JmV�鲉��œq�.Y�G�~�[��&���X�4��Qj_i<�~z�����֣�AK�}�V�V'�1%0���%�����c�l��[n_��n3�Tk�95ÝX��w�#etr)q�V�c�PԄ$��F��Y���t���T�)�p)�W���X1� �j/R�����`�ޘy���/�s�J^ZMx'߾��+�t�K!h�0;���}�J�u�G���C��Rk�Zi�Cf$�js4��ݭ�
 &Z=��qW]w;���A�r����HJO�Ѕd.�[�4$;��|��}��ry�>X�h�,r@��፰�W��1W�����`�vK�͢as�X�O$Dcz�eŹ�S�a���f
Y %sߵcj>��D�9�:\v\o�`��g���?/�TMQ�ѽ�<��<�תV���/b��wVzBc��V4<��a�2��^���WdBL�T�[mX͍�O�N��^O�D�⥪^/���G�F����zk0_/�Y�Yu˖kWD�rL�*#3v������n�\����z��O�#��S�Il-���s���'��\/M ��B9J��T��^s�n�d'��|�GaAI�M�c�6��SK�hl(g(�S��~nϯ݂u/l��iqP�fT҆l-Ci��tT.�b��~�%�{�mG1TVjK�s�����I�`&`���V��ko�kg1ۦ�}X i�-�,/kN��Ui$t�w��?;}�:�41?L��j�i4W:؇���R1�*��]�}fȨF6�@�'2|/����1��ؼ펃�h�%��@{�J��5�^A�ʪ������\��{RY4&a�Ƌrry&&��C��(��9�L�N���0m���7|}���V�u���U��b{7�ߣƨ,��yV4j��1qN�^�)����AS����@��mv �"�.��ʉ9%�&��y��E�ʣ�J�'�2V���0�-OF���%Ҭ�$���uؐ�5 R{�Z���h�פRȍ�����I"�d�>�s�,6ӶE����f�C���3�Qe�I��j��y�J;]ԧ��[U|���\����4|v�p�`{>��6[!�W�{���Qި�����]o����4���:���`~�}L�4��:�\��;d��n���;���P����q���`æ��?GG����wtI�k6%�!���\i,��g�d��*���cU���V��}u��z����H�X<�Ǐ�<컃(ò�s�~�|�}�4�I4�t��Ϊ�]v^���p(��}'�Q.d��i[�Sm�t��^;���n����\a�K�� ���i�ʩ�a�ci��RZ���mRs�Y8J�e_"`�t^϶�1� �^W�~w�,J�mo:���Ci���g�+�.�v�4�I��:�U���p����g��'�^���2.���fɰ���^�X�E�^�yG�*|�o��?��Ͻ�����~���z��O��gN�jm�@���p>V���.^����>z�n*.�KY8����?ހ��N��gq�qo�.si����S>�J��l&�~���Rd���7U�o� k_�(t���-�ㄌ)���+o¹�]�n�$�b>�c�z�;�(,�1����3��
������ ��b��Yd�%��"�nƞ���R;͙A�)������B��ʒN#�d��5�ю5hNgD����8`�?0����S�u��R?L�+5����*�������#�_�Q��������\h�����i9���L�����m�mE3=�*��ق��q��io�T^�D[B3-������+ ��a�%;�����ް��&G[�P_ʊk���0f���$3��d�E���i�1�>����dqs�v1ֶ��k�!4 kF��A!�gm�9?j���H�b�S1,k�k�S�|Zu4kSR1}ӫV��?&S�h��A>5��(@Pc"���V[��n~��"S\�4ͼRY�^F�b�[�^����,��k9Nz���cE"d5*1��g�k!vwLzX1P�x�h���{~~�m�u�B�%���T�~��h�#s:,�೙��ԣ#��Ђ����(��:̐z�f�<��&X�h'���J}_�	X����U+�v�1�i���&BJ�Vj\�B��y;0�D̬'�~����Lu��j�� Ӯ˃��<��K�c��� t���M26�����620�Fg���7
�WŽǢ�!qAu�Y�
���E��yL2[�S�$�Y�kT�������d�Ӑ6m�v�~��>�����/�(}Y�z�r6)��+�_��J�c� �_V��'��Ls$y5�V�{�-�#�?`�6�q�%<� zb#~�����밵�D�F��IK�A)�p��D���`s�Xe=��
�b�!8��@�3g�����v>0����gk-����<C��[_�J˓���jD-��c���3'�(�b�pC�-r�ϝ��g���8��X8��h����y,��_}�o���y�^'"��uo��)�vm��uՅ���?�ݲ���m���9Lc&>�6;�Y$�4D���5��\.�}A�A6�0�AlHg(M
$I��e:+2�>�d��PD�&H�"�2Y��i��&�V�;���^���h�n2b/zk57O�'�5*�Rv_�&U>�FfXAe��5�7<Bг]ء�����&ZS3�4[����P�<$T\jLI��щ�c���[]ј�f+�\	LS�����(O�v1��Ly��>��uM���$���5����o��ڍ��$qLL�J�-�BWމtu0ս!J��v���������] S>�W�rw��gN���F�����܍+�p/֮����FFG%���=i�!�Y���n�׮�3,i���2�L_V�~RUɩN*W(��O��a5��BӘ6Dc�<R��,H�G�=��|�����_9����k1=Ǌ��ǋ�s���c_�7�;F�[5�0���t��R2�yk�������a41�f/%USV}CA�m*����b͓���C&T��?�H3c��n��7H	�ib8�Yqa���.%�͢2
���6�|�
�'�J$ͳ��He��7�����D��]�~�Y����מ+q���+�0�����6.�����q�qG�mo8@�^"��SM�y���������=��~Fle����n�����~�X���Y��HS��·�/~�E}�[_���+�dv{����L�y�}X81�s�>;o7"�Q���Z���J�x�_�Jup��犰��頛ă���o|����&@5�J`��5��W�'F�K��l�;�7l���g7��Ě�U�cr�0%��L��!�I��:5�ʢߥ�)�����:M�U4>3�l9�p��E#aܕGD�z�z�E���-=�l����G8Q'���̰3��JP6�A)ӒVP���06T@!�>V��j�ƭ�eh;6���*�V��tk�.��n<�B��jm����vR�ɠ'��\m:�
0͠<>��TLMcj͢���?Ec�9P���\��4�63�#e��F�-��*#���43�.����4�l� P4�b��`(t�v��,�g�5��@��T錜�ZA����N��5�6�/��r�I��vA}V���^����s3q�r,(
�i�	�#Q�Y�;�W- ��D���w$F%����Z荴�ϰ���
�rw�8�U{�Oz#��D�&�q._� �J씑vVSKf_`fL/�\r�Zd�E��TV�t=׽�*�9��8�7��q�Z����!-��@ �]�+pIb]��:����4n���U�ª'�8��^�uD�5v@�����{��B2���?�n�/��_z���a��iY�L�^���}=H>�F�ׄ�F;�g#�
3��~׬�.=���L�$eZ����C�)S*hh�j��I�����&��[�a!EoT�1�3&� P�u���4�o��i8j��p(�c�x8���ð�6y�
����k�Bc��J�X%7�s-µ<>*�ٛ��,m����V=����;�Z7�f/�~f�l�tA�(�Y!	��N����2̲(WCk��ᘋ��H�Z��Y�8D̈^��1��
����4�t`�AF�N�WL�@4ԗ����bU@�����B\*�[ٓ�}�1��x��s<��$���H;7sm������}�z41���3���Db;�W0�i�,�y�,[G��DA�%u��T׈��,��7�4k5�*Sȣ��w^�v_��rF��t~����N��33��+e��@h�R���R����M���5X���Yג蓥)����!%g���dR����h:�p+r�����V������5+��w���W`�g>��47cV���,:���r	��SJb�E;t�U/�|�}L��7���|4?b�J�O��t���`����y�/�j�
lI�m�T�*�J�y1?�+�'y�JS����֋WL��)c�v�vE�鿜pN:�5��`ʊ�+����!;� �/�~D��ϐ�{� ����b,Sdv�ee��:��@�6�^��\���,^<��cb�R�715S���7c��B?]D���'/v�|���^ƅ�L�rR	�f'Q�^��b�x�|�4���49��L��͟������L�z;,�;O<
�9���n�V_\k���@6I��}��	��p����9��t��N"'�Hݖo��>�䯁����<�����U�?���Q�,��x`e���'��S`�"AC�R!�L����$�7!Kk�^��r���,�Z�_>�d�mi��d/�v����W_��}+����.(�[R�2��o����!u�ax籇���0��Oa�ړ����C8������*y6<d:�~z��p��`��W�� &F��FE���>��O`��W�k_9�ﶽ*f���~~��k�p�����Ď��H'z�8��.��F\u�uX0��O�M�J�AC7���]�3���z~
"�c������fC��:z@��B��A#H���覑�0�M�HZL�L�i1�jҵX�)"�wR��)t:�w�j@ˀHiX�<�M:H��5��>AtФ��	ЖMA��6�b��Z�Z�İ���>�J�sn0Y�o�͊�x��is@p�zosC i��H�M���YT{iTl������B['��	�r�5K��G0[���A�%����q�G�S�+�(Gg��A��^l8]Csv]�5�)z"�ώ�_`v���l�^�]s��!Ǡ��F{fIl�L��JG�uj ^R1 ���A��k��Y����HO8 B�S��a��h�B�����6�T��u�����u�F�!�B�U�Vj�4]b��p� x�̫���=Z��|�Ĉ0 Ĺ7� ��s��f��5�5g��^���=+�I�!٠��b�:,�+�z�#�=�	����m��G%�K�qR��&��|O`�H/���p��n���K]����r$��Sݯu?�PE_�OלUgl��܈P��IA�����yP��q��gL���*X��oh��ё�T@���b��#��r��u�:�C�Ց�=c{�r
�4O� E�ıҞ���qR�/�ou@)L�E�F#����Sx-cA1�'�LM�ip/&(�j.4i��S�0��<֩�@Z�.A�B����P�6+A�:ҽ:
��}�r��U�a��w��������y1P�6�'�8K�    IDAT�z,:b���S_��X��FS�=�y1*�O߸���|��z/_3��:�nq�gF>m$٫�R�wZ��/��k�No��Mb��X9=1u�D�,I�h��'1���fI�y�?��t�{bc�'Q�d�dX*�Mx(,<C1�Fµ�k�Y��i�aQ%�c��'�>�����n8z���X�|�4=WZ/�GR���4�d(n�����Q�?o\=g-�(;�<`*�$	�W�H&�����
����{�8>}��q�^c���/��5{����H0Ax6��2<Ә4�� w�m.��]x�M�w�H��jZ�ϩd�-������>�w��o�3�^�%�O]9�m��ű2�\�ɗ��4`�Ṽ2R�d�Qܰ��(1W��\"�<�>͏���R��O%���U�n�ƛ�WRR1���'�B��bX1mwМ�C�� J�x����iǀ��s��K.�D�I�f�M[�*������0��� S��$�d�U���������Z���Ӡ���,���W�cBI$�w�p!:�ʻ�
|����eS�A{��>s2Vn;$-"�7���W\�Wl����i^������ڳ[�h4�C^�^{��i�RL,F>�>]ԙ�Y���S�x��5�˝���\3�lq�`�|A6fV<�&K����Tg6��ڂ��q�wO�+�� +@ԿN&4C�g����3�w��f��˫�]w^����x��^���6����_�N~�5��3��P1+YM�=� x��O~��X?�DnhB6o� ��+��Xk�Ccz?���!��2˶�}��F���;�ꇓ>FG�U��.��4��)��Tf&�ϠYC�U�T�p9����8;o�C�L(����.��Z���OƧ>v� ?i��Ha��Ǖ����/xž{�3�8A+b�l�~rޯp��w������y�R�N���ƽ���v��}�q�yٰW�%{ŵ��G�� |��Ķ���"���x?���������=��~��g�\|����n��h���?�7�2+��?�?��x�iT�=�س}
V�t4�NN� V�Xg_άd��֛��\N*s�X���Y��I�S��b��B�(�N�f�)�SE�Y<��x�t��O1]���4Z"w�_$�*A��>�&��:�6� Xf��T̡TL�]�`j�zT���3ƄR�ײ��f�a�{�l$
՞&L�RitR4��&� 3�ɡ�H�kj1�m���7�[��5[A��tV*���<M�����a��)+���!dF��(f�P@����J�����6!���
0d��/w�Z�&��:�ż%�̍S���N� 5t^�
��#K�FﴶF޻�!�1*��P�x����շ`ߗ-�WO���Є����0��fc5����֩%[�3p1z�!�ΚLg$+K����R��	��v�n;�8��"�ƯA�yA��m
&tl����3x)xl�V
��!ѰH�<O�=����ŹzNӵ��a�tL�c����v��I�QH!��(Q���g��Fuy4�c�����+1�`@���`l���AZ-���g
�Ad$'�T�%�4Hչ��'T<�<�,��|������O�������F�Ǚ��8��R���W��~�V�4��Ii�,0V�mj�.�hǪ����`��+�����~�g�Y(�h��(�r�q����9�s��K�=�A;��K����l��\"����p�+V�5����Āܒ="��[��G6�	Zɑ�H�N*)��Wfk�]��g��_�x�<�yz�V��yt��KQg�3-^Z� )��SX�A�����T�)��WRڊ�����	�NP�qO�#�(`�Y9ֳ���������h��x������a�'|�/���+��~i���}�M&׽*č�ޣ��<�����-Qb,L]B&�޿�Nc��
���O�l��5�3A��%]bTp��'>��i;wᖽª���)܄1�ow�kV�n\����_�eEō���5kU�~���/[.��ޙ�&^aU� ?��wϹz��8�+"I_��D��a��
��:�d@`A2��Ma^�x��O�J�=d�i��:N19ˤ�,�<('���c^�\����n�����zS�	�2�c?T`9�r(��;L[��V�EcZF�T@`S��R15/Vl�I�5��o�W`���r��
0큄
��k2P�����%�buel ՚��L�|¡���`�����[�	�&uz5�?��s\}�ȤS8��pڧO�n۔�A��$�\v�]��vQ.�ϱb��-(#��+�����#{9&Fu�xvHL촻�?s�\��������Q撚.#���4#��l:--*�[Q�Z'�bvX��9g��}�meu����ܙ7����b��
�%`GQQQ,��KbK4E���h���%*FS�K46�
�%D�*<�+�n���Z{���`^^��{�9������k��׸��V0��s��~&.���X]����G�W��i8��㱅n�3���n��8KU<&��>������Py񋞏Ù	j�/�+W�'���5Pj,�X�0Q3u�nڭ�%�T���3��hX�H7g^mT��3n,.�dD"�H�h�r~ �r��l�ei��`�Y��a�Y�|�̖���1^��S��O��vn�zw��}�[q�W�%�|���K�	��{ׁ���Wp��~��۷�9�z�9�n�p�J��׷�_����������?�ر�zTo۳�/|�\\q�5�'8�����O| Z����<��2d���?{�㰃�)XQ���^����1��9�Q'��/x2Zu������?���t���g��;�HȵG���?�g��}e�.�6%��a����@c����LS!U�������嚁��d&@�?P?i�s�Xs�h���|�z]�=��1��@O׀��P�M=.��fN�4�s�rT�q�9M�̥W�W�01`:`0�DW��tV���F�&Gb��o���5�	���f�V��J�����q���F�lIC�g�&��w����q���qk~/ˡ��E3�C�ֻ�;0�[^k��p`�({�%u�ꔀ+ꔷ�0���-�M;�+]iq�-����X��K���Y`�Ny<E�?���iN�����2��I�j�9�r´-L�Y�&��c_�[����)c.qH'���k��QUa2����R�=�8��#�s�<Z4v��M}�V!�D�C�-Q0�ê��Oq��.��i������'W�6��:��L\�j5���AC:&��T�=<�w�iO:��Z��^��\z��X@ؓ�pKu`<�̰Ҟ���|�K�� ���pLL��pW欟���ʙ�`�6�V��m612\fY�d��R���d�6N�{����>��瞤eD��I�r?Z�%���o��1���\�0�T�v��thzl�>�  Rg�r���,�jii��ǆ�߮�K�k(�5wNh��P�泣�P�kT@�S)�C�gpõH���Ba�}ƸQ��N1�j�+~�6Z�}��]����\���{K��4�Ԟ��|�\��*`�\�l�"�[�RDkIs�v�,��y�t�>�>�Ľ�u�8�@�ܺ�m[�4�4�t�FL���_�<���x��[��ֽ+�Օ��=���U����m����OʘVZ�O��ɾ;�<#G���5��+�ל� �!s6S7-x���jt@�o�ۋ ȁ!O|T��=�;Ҍ�u��uB<?#j�c��)`�+W���y`j����+�"~�Mu�i��P�$29�V��Ŏ���c�,|ܱjj&mQ�4)eĶ��ތ���V �����2�~�U򢓬g���OIʐP1�\M��D}d��S������]�B��5� +��C{++��ۘ����> /{�cq�Ί�������ȫ7�y�M�[þ/h�u������|���)�}����o�c��F�c��h�z���S�{���h:Y�s"�V�Y�^o�"����E�,4$��m��i�Y�]��g��z�ָ�;�T�90-�Pٲ�����I�͕��_k2�'Go��G�L���b�Z =e'!�%Jy�vnۋa�+��Q3-��T1,L|����B����l-����3�t�5P���8/x��L7U�7�W�1e�/`�Og㿾}�FL���+_��;0�T�������%XYan��j�����C�v����>w9���c�,���\a[��!P���|�+��W��!:����1fOg���2j����Eg�V��{%A0=� =T>�kn��-��0�w��f��1�w^��'��'=@� ���u�����3�}�}p��N��?^�=|����O^�Ǹ�=�.&0��o�x�_����(�Q�����FB�I���b����PM���J�����J��kx���zJd,ѱ>%c3#(�R�Y.b��_�	V������[8���ra�Ҵ�Cv���m44)���8
{�-㿿��mw����׾h�v��˯^�G����U�U���C�Qw;[��TI����//��*�s�먻����0�����o��-��,����bǶ�q����G��3���p���E�{&����`���O�����s/Bw8���w��صc���O~~~��+��
Nx�p�c�R�B�;�7Ͽ������9�U�9Дk��T������%6�Adߦ�n, ��R6;ڝ�=7�,-�P�Z�V1?7'	,���NS�}}E��ߨ�}!��+��Uy��U5�Ӻ����A-����>�}:�xU����5a�z��f��J��[o�U�m5J�(��!�f��w�T��A�66�4��0�Dm��l`��z��1�r.V��8���wea>��T�`*�8�� ��A��_�a�n���\�r=��\�C}���ES1�ѣG�֔��-'�LP�1�}:��g�2��=z�?��i��I���ǘ������W��h����z\���=�>h}�:H���������)vlma�-ZW�Ş�|���j�#JT���R
����.�d��<�l�� �'K�e��Y��c׎9l_���\�G�#�a�)��n��%m};J&3���p�շa�� ���h�/J��Ā�|��H�rc5(�Lջ�kJ�fO*,Vf}{�ᵧc�:I-V'������g�n~_��gFD&�Pl�7�3����LB��[_VȪ���z�����Dy�'s��a;�v������]�P9���`�+���D٪6<rR,�
e��"��UQ@�	��Y����yz�I��@]g�K��:� ��O��Kg�9h�IV$����Ҥ����u]E�#~���$"!?�Ӂ�d�ꩇ��WK���Nr��i��4�c�[&�G���q��;p����QG�#=K�y,���8�+�&ۤ�\Xo�������a��:n�}�_y=~}��}����[�qG�q�{�h�_�����s�R�.r2F�zQY�u�^Ϫꌱ"�Go����%�������s{�B�T��P�P�㶊M�J��*�vs�a�h+H��c����LS{������ �����
��ogAPAsD79$�� �d�q=	t�ȧ���R&�1q��`ѯ�_ǀ��4���㛈�(eF��=t�3�1`��;�#<���>�Ѹ��5��	NF_o����)C�
������_f�e�-IM�����ek8�?���^��B��?puS�(�P���2��X��m�u�{��e z��h��(3L���V8�T�f��Dr
�3��	��6F����u!�L'�"g�F�����v�����诵��٣�q5wL5g�땹�̓J@����{��9y~ՅfՊ*���R�d�
�Vp0S�_&�0�v�����>�x�k���w~_;�G�R�t�}�/�:h^7��=�L�/}�b�[�`q����|�N��N;nuÓ��[ۙ�#؝`p��:9v�������|��f��z�:�2�������U1%0=�=��}�+�ko���g��]�յ�Z�s�C񊗜�'<��3���K�����2�~��㤓N��s���[���|�?��8����z .�M/݇��]�9@�1���~b�����`J,R��"H�i�=��e��e�������QU�!���}�X"h�� /���Z;vlS	}y߲�K�L:�1�dw��Њ��q����l�0���tĴ�jx�I��{u��9.��/q�/�h�^0��'�R� ]�?��L�ٴ�=jsRc�C�A�7����2?�4v C��\���q0�}�#�s�4�sX^��_:k�)��b�����	�S�+�d���4�P���6f�y9(��|<�UO%�RGR&�L(��56ՇCr�͏f�-��P�Ge9IW|<�x_գ�RTKm~h,g��ݎ;XaVXU5�Jr)���Y3چ���&C#J�p)y�H�	��h�:���F��@�McL�V�l�]K�9���0�b�@�����,�ld�����R@�R��%�@��Ot�v�J;v�ƾ���?�(��-`�须l���p���j����i��a�ܓV	3�]q�T�[2���H}��6tvfF;��j����J�?O=�����K���g��HB�����4��}�|��e��Yۏ�k�-����u�r*���x���ѽ?Sc�j�H)K�͞N�'#Q���8�%��lL�F���~f��\ї��A��n���3ޭ*�f풅�j��1FK�Y��*N`��j}�z�ܐ�ɱ�$�HY,��[=�4���gJ�2%K4����p�4,�L�$!R�p��`OTE����`o��*��� &5F)�u�gJb���r���<��Xv	�f=��bf�O$Jί@ױ��ż,��Wkboƿ��&"#�$j��f�DR�J][��9I�vl"~]I-��j@�_�+N(��CTnĺ��{�X{"i��%�2��l��'W8��^�*R��W���ȍ���gYWRE��01�~Me�L�A�Zs�_�kbi��-[t��\�~�k�Q�߿��v���`��ۈsQ���7��R��5�Z��P��\�ȳ�jch���]{:;�4��w�e�уM�:�b��&6�L�ƈѧ�r�Fu%ࣀ�k���I�l����*Ŷ���4oD����U��E=��syW�<`�}m��e�A%B#���L��Jo,� �YV��'�k�]�;�$�w@m�\��!W��}A�6+~D_�q�Zf����z4L���g��Y6�L�,Op�R's�����ȝPeO��j��6��6�Cr�'�t�]�f�:s�m�<��K�M�_���O��U&���α�dqK�DJzvdmV�����AB�:s���H�XŔ��%��4��*L�/8�7�J��u��Q1uW�b��⼍Ǔ+/+�2>�&���Je�1ݿ�b����	�N=WRyx�L�L�r��r	��9���^ň�.9��l�fԇ���TmMF����8�ӧ�b�@=��0�ݦ��|������'�׾��	�^;��<���h�{��O�k{�y�c�̧<,?$�tƹ9Lm�}5qq2�R���A����3_��Q�b�Z�jY}��{~��x?�v�<>�����mS>���c��3q�E��Z����Qw݉W��4<����"	J;GS!^c�Z�p�-��s���=��8tׂ6H����>������P�mQŔ�+k��*$��(�:3ne�Dɥ���P6)�<�}�z���Q��%n\P���BG���b�'N���v�؊�p(`:�C���$R>:�Q.	&b����
�em��|�x"�$^�`4��z[��fK-�4���{l�Q���  '����XREORK�
�_�j&�U�&j�g����8�Q�U8�Ψ��o:��g���|�Ь7sf�?�Y,Q�K�!`#[LB0� ����ՍG4~ī���V������a.�%_����)��9>3�|t�"n|a�S]Q�G���L]�;GΩ>��dy(+r\��^/ę,�%#f 2���<Z��N�=��w�r��,���2�k�[#(�k�];A�0Jy��5Է-�F�ԁ@��r9Ϙ�
��`$�9��b�)]{U1�SUޔT��ϴP    IDAT�}���C'L{�/�E�m	�fͤ��g9����?\�#kh�D3 ��{�*��%�3�4�ā�D	��z����NYI)��F;�%T9v\����-[�P���%uL�C�=�m�r6�h(�mՊWz�*C̭�o��dy.�+�Fʛu����X!ҳ��K����Ýk��G���`8��ND �Q~/�L L2TŲ���\\�w��G�>'s0�Mk=�6�=�{N�'L3��=M���^��Q��U�Z�bX���T������ll_Erb�\���Lb墩��U-7��b�Na�!˫]���S�8���130�L^]` IĚ�?	��B�D|�F0�y��MK*,���8��>�8W�ؐ�{��^O� ȥѥҊ-.�S�k�_�#�Ԫ�v��S�}�{�J'�+��>��JB$�|]s�&�kn�">\��zײ׈��b�߀��"���=O�3>�D�+K��^�g��GN1�	���w��a�+�ʽ>֬je5�y��uL�RU�gq�DҒI6[.�V��Rl����mj��x�Yu8������� n���OME��H!ӫ�Y @�c(�z��ދM��2j�iE�;{�3����{�}����	�ͮՒ�9�y��;��vAJ��1���ڳ?����J���m��ukW?���PK8��y��n��JDPT�rj��_��X ܨf������ҡ�˼�7$��(��g�& puG�9Ҿp�1�3��5��>t��p�]J�Z���|{�x�:n�}ñ�m�7��گ����Z<ۘs�xa~����Ԫ��}�|~�bY��c���u9>�o_�`��Yi�9��!ck۔tvv{/�ǵhOP|��[�BD�ݿ���s׌y&� nͣ4�T�3�i��1pG��P�Gm�����	�Z�t��9�a���0��LEH�՗~���y��hs�đϟN�����~�^�z}�Ƭ�ڨ�2��Y�Z�~N��+m��rƺb�6�bz`��W=�DS�fX����+���H��g���������1xݟ���d� �p;p�G��/��w5v�<Y�ӟ�p��e�����niv��騰����m%���p+�O��8.��Mhkh-n�F�.cu�M(��㮇5���n0�~/�wo�.��*tz�.p��x��'=��8lgMw�	�E�gػ���}��8���mu]�2{����9���>J�E��*`�r��n� ��x��6�@���I��6^%�q��f��f�.V1�Ry(�C�w;���Ձ��6�	�<p��+�k���uz^��$�4I)DV�T�B�ՊY�*s(��t	T�-�*9�$A	5��|Y������Ǚ���f2�q����V���
����@ŠX��u8�VnJ��Mjq�A�3�2��J6����Kl�bO������x��	L晼�n�A�`g�����ԛQ�0���r��1 5��r����IB镠0҈ꗞ�c��|B����"f��'�5�m���C��R����9����	���(Q�)����E
�(Β["�A�X�3dŔ}�f�%���F���R#����Q��[YCo�*��۶0Ճ��PtY�Ú[� ?LI�0�R�[ݲ��|]Sِ�:�*)�^1-F]$��eʅL���b�bP~v_V�Q!�X��nꑅXc��>�$�Y�ϫ�NFX~󐭨��^�b8zh`,����+p��%���� �"Xm7��EiVL�,��mgKr+�����=�u��/��Ӏ�Ԩ�X�I��gHY���I&��r�9txP�9_��o�~D�HH-�	`B`1V�=ey��Qo�e�r������l��H)W1�;/��FM9_�C���HAk2�;��f1� g��4�u ;�m��?s?K,7������aT�3%�`OY/Ԇ1�Pi�ǭ�O���FJ�$��E�^O�D�����A��m�z�p0	(X=�Q�/|=S7H��{��y�̱��J�3 ��Iҭz�~'U-g�VY��ٷmD��c�]�d�N���;��5͏���
G����ͨ'\�-��ci>%�fB�~e�v��ʌW4k�خ*2ך�q<�to�_T��N~'ii��6x�E��[�^�z�I��~��N��l IL.�g��'�E�ϑӰ�e��:j̣Xf_9?<���Wv�r�Pmv����S���<���_)?���#UL����G�80��w�zn�'�{򄈻�Kis�����M��z636k"n#'�_�Vo�8�Ǡ��������$�}N�����3K�,H����~ Sou����1���q;�S<��Ƌ��@�4@b1�*&�~����~��n�F�E�%�!���L����&Z��^/���4^��/��,�*#?�뢀߮/��
g��(���8�\�`2��2�+����p�͈�XDR�H[��)�M�-�1e�q��SUQULp�ӄ�9�+k�ļzI�[�ӕ�昚�d��Mo��5a����3�W5ŀ�ql}2)1U���3!~A~ �ժ�qG������y���%�i�¡i�9���_��'Π������(��5�H<��P�������{ӚUL����	�|�1��W>��l�_}��ؗ��o]�^g;���7�'?��4��#|�,��eI��Uc⦚D��#�����ƻ��\������`���2��܈�d�v���S��n������%z���XX(�~���9�~�q�#v��f��f2��ؓ�K��ɏ=	���	�^��K��_�!V����B��P�C�\$MZ�~<[b�N�t��(ŋ�?&�2f�fe�Y�a��@��7o��Ts2�`8B��ŀS�N�hs���<`�����u���	 QF�#����^dX���(�t�X���=(���Y[|K&��z8�C�fR<�%%��@�u-��&�����J:�Lo2J(���LE0C��C�!�:��K}N��^�w62Ώ��p�"�dժsvύ9f���!�QؐnY��Y�6!e��z�덦�s��v{t�Ӊ����gm�=��I�3q֍յ�9w�J=��`��2g��� ���~��!������)Օ��=1}�j27.�d̤��L�S���Ȳ�ϣ�u��U-�n��mk�sH���	
4�ZYG�+I)+���&��JN��'�z������˒���޵�w ��y�s`��e9`J��`���n9��Y�N>�!W15`��-�*�����X�gA��J�Td�G�|�/1ў�8�8ST�i���7H˱�QSf�^��Fd,]�grYGt3c�cf��P��n\\�fo���X��'9�s[�DJL�TB�9�$���EP9W�7Dw�#%�L�&$LL��ـ���n ����ò>7>�pbo}�D?�)�3 o�X��P��CW��c��][X Y襸TQ��ek��ݒ�̵q0���^�z���Ŝ�-
����<K�Ӏ����fs��0�$�e�%��2θj�C�?�t��0��/k�w��+9��*�~;sD@�U�ֿW?s&:"��P_����|ܓ�{��(�*�7Y�@P��K]>"e�f�hF�;y�fgcH�3����'��y�����%��,��H#"M�(3�۱��Ώt��4uٱjS>O�n6#�.��C��*Cђ���X�6+>gg�����I�U$��jS�0�B���j�!��‭U�刃Po4p˾e�޻���)���%#�y�pѩ�|L�%�o�)PF�D�ҫ��<'��7>�{>��$=j�wگ?oRc����c�G�=j�߲����Hg��-{F�/�ܐ[�~I�Im� 6 ����*�f'�x|o��fʱ�\����U��}�b���K7_� �#A��1�����}�qx�S�Î*%��rQ0Y�����w�����C&S�&�m����S+��Ɣ�A�U�(��2{՟</}��5��T�SL
3�Q����7}��э��Pk͡U�O�Y�z4ɤ����d̢��ɜ=S7?��Bk��r<��_D��=�S�jI��0\]ð׷$�J`:/p)`�62{� ����ñ&tW�,ׯY�)n�jI�6�0mm�k�ZT?1�b�)ߟR�9��9���K�d~��.R/k�rD��0Ÿ�����^��0�_����tF�����߾��{ᥨ��8�a�0=t{]��W�p�G�����!:��8�G���|�Q�gS|YBK@�����v�Ǧ%P$�v�
�����o\�T�D�7Fwu��w�Jy��������.-<����G���@�_�h���|	��vm�����#<���0���l��������n؍�?�9صԢ�W������|�n����I�f�r��\7beakS`��ȃq��B	o�^�\�8��
���Є��Bt�{�b���[�%��	LW���Sp���0a%���ɹk�K��r<f���Z�.��h8BaB0dUN�&T���[�~��y�K\�Nn������$�9i�ƺq
�f�����'ʈ���zgB�A��:$7v`%	_P���f}�&�5����<��*�m��/C����|��`(5GȰד���O>�.�qZ��v�Y���fdˣ/�B��*?[\�=7�WFU5����s�&�$�-�0�"0m굗��b�11v80	K�Э�Nd&�CL�Xoh��s��ɘ����j�S�N��i��dpn�v���4�r@U$g()�3�����PaC�b��E�#P�{�uB[�Br�%0-<�8���Qk�i�r\���w��ڗ��>!
��Jc&�K�.�Y��9f�#� �a�z)��*�g��`��Y�}�Ϋ�'�o�&��9�f���p�ʙց([f.E@ĝ?*1�}��=S�L�Sa��N��zx����'�����A�,�9��[�J��ZR�o$�q��6%��8�N^���7���ӓj�i>qV�������w�_�Al���l]��(ox��SJ�8�P�G�[�A�^�P:B]Rng�͕��&�^������Y�W�=����jcyiH�-��Js^�gy8��k��� 9��q%κ$��.4)��`>)��I2�0�Yz�T�+���q2�Ԁ⸋][�8|�6�ڹW_s=vߺ�����92�n�%��w �{m��`NZ$�����2�䠖�?UE�����p紽��^T��z�[��U ���$Fm��P����;�׌ͳ�����V�6�xN:KmE�D�sp'^I���3gs�}w��~l�p҉��3��H|`Sߴ�g�6��g8�GWcP���;��Z{�@���Q�Φ<2��XQ��^�P�@��,�˱W3�l^n������\�C���wU��"O>m�S��2�ߞ���P�eG���<ynW��E��_מkƊq���+����O���Qe6�.�W���з���T����tј���N9/;��^��3#�FӢz?�������2��e����s$�S�#��`�U%�~��@��fu��B���E�ӛ_��{IF5�E��E�π�y�9���W�?�GkiIRU:�F�0b������P�ԉh�4{ץv�OtX�+/ǵ�b:��s�X0>�����t��B���TU�(/�4�@�����&���Ű�ʁ)͏�V�K��!��T:�0My�7��ӊ�����RU�g�ǌR^�A��x�L���ۙ1A=��5�(�bj���fQ�{t<��s����L*I�)�����%���]��g�w��ϫ^�t������b�����U�|p}�,��z��~��[�u�ŷ��n�;E�W�����v��}��aM|�=���L�����G?���%�۷5p�{��=�^x܉�a�6�8��=G|8���r�z�<����j������x�Y�Ï�\ư�����M�8eZ��brX���S����|c9����<�_�k��R#�K��Q ����U��u����-�K�b�{��fhFE"�^�K����H�#�x�Ix@R�KWې{�F3{UihD"B1�H&K%��ت��}N&�e���WL���_V�-	#h-��ki뢱��)������5z��
��G�5�U��y#"���j��@-1�X'��f�[�YM���M$%��� K��I���/N��gR�Q(q[�����~��f��o��ĉ$`�c@�J}Ƃ#��=�Oc&/�)_{u�*zڑ�����%�Z�^�P���8����G�,��_�6�:u)G���7Lg��b�"�eR���B���{Vό,�@-Pw)/e�L�^��-(4k���3�)�Q�T��K���-�Qt��UL3`j�����gn�"�S�-��]F��/O�R?���b_�_��\WPk]
tJi�{J�VzT*��k�8�)0�H��,�=��w��J-^9�1ZN��1l���d��#JJh,m��ZĬbR�����m�~�Q�B�7ƨ�Ä}+L����W6K��b�p�����2��ң0UUѫ�[,��$0���Ѻs�.��U�\^�^��y���F1"Z��p3PI�!H�\�,?JTLU��K�F�N=���I���b�U&�3n��l�רȥk��̊v��R*NЛ�y����S�0���=�C�z�'b�����κz���%*��
{1Y��bH��s�!�w�x���{��s �&qU������_�ƨ�Y�t��[�9�k:p��m��8�{��y��!���E�v�A�v��̂�ֹ����P���eČ��8��B�����|��ѹ��X�y�W�&"
�2>�)�,��8��F�ƫ�>?�3� ��ُ��K@�vV���K~5�߽�SX50��R�lq��"�C����@Qv��9���N��}���I �*��Z�ui���{��S9�<��N�=�@_�9"����"U��GӾR)���3o�!�����0ȭ���c��:�i�}��^jҷO}��%�
M����nB/�U,�x���˞�p쨳bJO��q��o}�G�o��-��9�si:�g*8�j;��$�ֲ����dyy/VWn�����^�՟���=��h� �����S��o?_����csh,,�얜7��{�s�s�QI�:�6��=���3`ZDinNf�c��̑r���t�15����c��&���xȃ�--U=5KT�Y��YŔjG�1_*'��ɕ���#.��5+���A���	� ط�S��@�_�wT��m3D��K�/i�H�6��$4{LG��N`�����Oy��>.f2k�፫���!�{��ШW�������sp�V��^vMg}�s8�܋�~������ 5��X&��&�B8�;#h�Ǉ�c$�|�3��}�?�����������c4\C�������{��K`z������O~vݎżv�<���p����Si��O ɝ�\�Ȅ��x�|�[��ß�.��u��u��%'�H��$W�s�0$�bǃyW��j��F���' �t{2"03f��|�~V�tڳ�M̑rg�ެ��l����x�,���E��TO��f��!�I��z�n E�ʒ}�Ȑ�a���28�i۔V�2W4[�!����	Wf��j���̉�z��-l��Z�L4����)+p�CT*��*��<!�I� �cX�gK��O)_�ˎ!�|�9�e��_3�]�9�F�761z�=��/�*�Y��Uzy��_b2=O� \R��ÝE�>ʨ���Z���bã��{��v�9t6��"0e�+���g�ƀK�-%��=�-�˰�$���]TUt�kg�H�t!��r~O(�0`:E��n�ն$ΥJ�m;P[h����>�&)�tV)E�9�=M�)�,�roڸ3?2����-��x�����%�,+7�̏<�� ���u�bDFR�[Ϭ��%�������`H7s�l�\��7f��������:��L�fr� C\Ȅ���4h2?g�'ڕ_&��}M�r'`�`-q�FB��FY� 5�#��A�ۖPhV1��E�6�5��fJ�\'��o�7Ơ��L�|-.�i$R������תq$�
YPI�]e^Y"U±պ��|R%�M`|�����F���­��Z�� ��p5�X�pn�F�o�M���9ƿ'�~$���se.��l�Y��p�4��,F�s��D��s&�sB9����V�v�(^M    IDAT/$o���Q�+n�.x#+�ϛH�t䁄�>�E~�#u���0�XlJk<��=X�A���KN�#��a�)�x� ��	��}���tf�5�P���J��p�W�C���ĖV�,�Y$� ����n��c��<� ���<����rʱ�gO�����4M�s,��18��M��T����:��%(C"f�Gwm��=h����=��Oy���{a��9oR���2,�w�����ݟƾ~]�TS����_(�ȝPl$`�{.�לbXNy_3b*�YE�����=<Gd���|�1:�f}q��6�Oz9"C��$W�������p�Y�����cvN*�c�����WE�ſz�<���̷�����9z�6�h�t�7�A��m�ﰿ�-�.���Ë�q"v4ITе�gv	��2���ø�7�(�Ĭ� ��]��ۯ�ktt�:1c-?/UE|ăQk�������M��g?��bk���� i������ �h.,���(?��D|�P����3�Pz�>m$�j�VS�t���Mu�����٪��5�x�\B���H��kw�.��Ң���
{T͑�c�4���p�!������u�1�	�tF/�rA�7n�>_��BV1%0U�i���JI�b�$��Q���bK�]=%������+�Qi0}��Zgڝ�W 0���Y1�� 1@ο���.E�VƓw^��g㐥���~��5��o_�w��&]|��o�#��zq�>�M��Ǧõ�-ѷΪRQ�+�0���'>�3|��`��1V��ǰ��J����ę�y�s���	���gᢋ�D�7A�4�=�: /{�S����Ҷ�6;zB}�kU^{h�g-����YܴL�ML�|�=��63wA��%:t���S��-�"��4U)d)aee�+k<�IY.z>��V�`n��g�X��L�6���P�����JՓ��O���D�o,i��*D�8T�s�4���o��.����mf�R�&V�2'���[:��G���Z�QE�H	��[��3���p��z�^?��1Y�r��!J���%~����䈜U��(��k	��,������M�~�أgE2 ������0�A}Q!MJ.����l�F��#�g��4�ā�'w�
2�b�3�2,_O���׍zLg,��/`j����S'7VVL�kX��i�iQ}��s����_� �xP&H9J����F݁zL��@�R�jIR��d���_�-���V�0�$/��ZM`�����j�d�4N�=f�1`Z�LӾ��pDaM��c�	��*G^?]�e������B�o?�R��d�>N2s�]� �}%0a�|�+�ٿ�w��2�_�ڪbe�r���R���wSZ�^�*?���MR1����%�K���E9Q3~��'��Ox�Jsu�d�kftg�A��)����XϏ�2t<�3�����"�X����k��m��%�Y�IՒ=��D3vW��n�~�S����`��>|	;��'�~�J��6ɐ�>�eU,/��wr6��VO�5a0���L�F-A2����3Y��l�w���zr$_�j��該%�H<+ϡ�������w� t>����` @q��[#W=J�2zK
M�*���^�ug�y�sp��\9�s�������c�맾�s/�RҾi�a��jU�{���C�NF���NNy��;�{��jp=����̈a�����Mw����5iO��@{�<�y�1'ߍ�d z�\��z3-�$7
�
p뽥�Y)m��Gom0؏��k�䅧������`q�����o^��}�|t�[0�LU�,��ѓB���|���eR��1�Q_O�Uyk�Eܴ�~z9�odVVyΈH[�Q�����IN��}��%6ZZ�9�Ȏ�;��T���d�GT���:.�g<M�2�����R��ٲ�HM��ɑ�UL���5��ʨL�[�l6������!�{��§>�\V�b�7�Gx�?��ko�aRފI��Y�T'Ҝ��i�c�����5μV���
���]�����-x���׽��ٴ����E�L��z˧��\�~��Җ�)	W��\e�@$h(C,�����ko��Ѻ5�G�Y*��:+�4����Gf�~$��������C��W4g~4��b����N9U楌#�_~N�0?���]]��P���В��O�"���D���.��r\]yY1m\Lȝ#������O`:���Iy����9�N�Tŭ'N���d6��g�R�7�b����|,^��g�7��˫Vq��>���C��c���7��+*^ ��G6y!�mq�r�=�a���7����/܍w���ؿ<���{+���r�=㽯��~o�?���������L�;2���� <�Y���O<�x|�cq���Y[r�c��`�����	\y�:��I4ÔRB;���o��2�.�|�`�����5����z�d_YYÞ��4S�I��p��.弻�8��\�l�t�e���=M��^Ը�S�؀�4~��P��Zi&��7YavϪ��&X���Ϟ�����R�����m2����ཟL���k�?g34�ule5�����1�k��$k�/,�f��L�۸���5?A�����d�dIF��9V�g��iԥf���%����K]kUU��J�u�J`��~�Ee����Q��+�v��a)p�
�u�� 2s3+�a��j�+�t���t�]�(�Y0�����h S�Q����sM�i~T+�`0%p��[� �N�S|���l��P�H��ގB�,c���ˤ�B=�����h����ϪL��[�����tӜ�A�*�r�+���ﶀ)͏t�q\m��(��F7��:բ�u��E�F��fJ��Pzv뿶$2��H�@2H���`C���>Qw�V�ܐk�]m�l5������s֧I���X�H�ߐ!��R�^:�i�����}MYmr
$��a�^�R�I=�FrX����x�\�t!$��NіY��#��p=���Hՙ �� ��a>�S��g����h�8���󊙪��?L"gK������b�g�6���%E��9F)R�u�u���z�3`	N�s�o��t�e��}l��ث��@k�g�;���1ٸ$�Q)�W,7�S=�MU�|���t�	+;�\��$���A麕���dcB�˞Hܯ v�U�T�1�W�*}L����9Fr�c�0\�!KS��/_��*���T�)ОW�|�K��}	�5�	+TUj��U�2g.3�v�"�]Ĭ_c�j�k�~C��fZD�`�֩�6�Rr����?l��8���~@�Q)湢uĬ@����ų�2C�j�����
\��,X��=C��l�v��h/��q���ƿ�#��qb���c댼EA#�.�x�G��\��^�r*�x��)-���=�����۴��LL���}'Հ�#}r&�/^s�9�Z/d{9�8�GK�.d��#��@�S>O�"R~�9��2ɪt����ʑB�P�*��i�T�<0��j��T�r�w��F,�+��%ŭ �.���P~JTA-�l��R��=�x�S����1�c���C�û?��o/�7��Uy�p���-)�&�|�|QH��L�ė��"��+�w�oQ�ݎ��t^��g�EVu'�~B)�k�����E�a�E��s��ڟ*L��u���9�L����7ۻ~ğYd+�Nk[Z2ҸkW�Y�g^������������{DT1�T
�x�j��N#<l�i�+�t��s<�V���G��.���ŌpLO=��>Vn��NO�fxΗ9�\İ�q11k��V��]�o�g��0�b���Ɵ=��x�S���wb�D��f4��ͫ��F`�K�5k8��c񪗞��VR�ŕ��ȿ}\�4*S�����c�>e
l`ۭC,���I��.�.$s�c��R�����[��Yܶg��}+�WQ�*�vļ����on����A����h\F�V��-U���#�= ��<`	�j�j��:P�&vc��	����}�S\��5���o�ڛWQjp�p^�9xF��)��D$~�ĭN��t���O3T���rz����������J��@MlP�P)�){j���1ѕ(I_|�H���6�1��2�d��ܾ��`� ��j���-� �9 ��fx�m����O��E5��=�4Z[YǨ;��ɀ)?W�����e�b[��"U��-O'J�E5�
3�o�r�v���
F�0n�*�%�����j��*)M0��p�xv�<1�����=%�o,�����������BƠj���b&�i-�ə�?��b�����)o��[�V�*����ܬ�c�o3��mQ�eŔ�\"x�h�T�V���п�Q�\yk�֣H2H� I�3�����pm]���I�df K-Le�h��ۭ%��#���r����4O���e�%#@;��|i3?gc�+E�.ޘ�{U>%�!��)4����@��\ʫu]��K�FC�nu5CTD�"� FC�ؼ��K(R�)���(VJr�\8�N-,nѡ�J�	�������b/Y�s���v���H��=W)ˑW3MijW.�(1ɧ�p��#qD�n'g�U�.3�)s,��o�s�%w>N�W�%sJ��k��+`��{�G�wW�^� J�����Ff��d�c��B�2p .��U@0��ꉭ�sY!$���R���׌�p�b{�	�&�'�#].�#�����<��6II��|��E�4�+9��d`�H���Y��XM���S�|�4��$�T��bB0��I���c4�_�Wd�m�YXé��/���bW3f(��XY����� ���O����5L���U4�0�Z�1ge�*�FL��%�O�Y�u%VC�s��D �c](.��'fcF�O w�EsV9s僟�FĚ�?W ���S��F��\EȸQ)$GѵWW�[[Ŵ����'w7<��ĉ��y�/%����PU��6����W��3��@Ֆ�o�T'�|Đ��=v��k"�~ R.�������ޛhk�\��?�� й���'�����(Dl�$�W��!�B��'�h
l���d��;�e����봯[�2˒[�A)��΅�,��@*�,��lc�9�3�M��c�D#l<�x:ftѧ����z���a�և���]��������	F�E+�(k,��a7s�*<g����j�WͦXYً�����m8�a��߾�8t[A�D��Ê�k��q|�����t~��}$�]s�����f��0��c�H�XK�F�s�^���vT�ө�J��Әa�R�|�$����Z_8z�ఴ�Be��q����}�F*1W���su8ByU�T����j�K}��T	^���E?�z���0�����V��Y@(�90-�|2�Ό�љ�t��1��Yw;j]��Y'�߀�h�eT0}�[?������,^�ga{��ف_^���?�9��P)���>�U5L�fj /�M��w�B�-�qCۆ1�ww
\p�-x��$`��g�#2 +8��>������Օ�w�������ɥ7a<�P��jy��h�Y��:�-5Q�w���x�k^%���Q����{�K��eW\��޼�koZ��Y���S���%?Q!	��F�X ���$�7J�y��ƃg���|���D)o�fC!}��rY�f�.]�Th?dLi� ��6S U�����"��#\���f��9��v�6���-8��\�����[�i���z���2Ts�$0ݲuQ�K�&��v8x<F�����ML#���[�r���IJv��%���D�˳'�3%�6�T�D�2�#Xn�g
���\����q�Ⳡ��c�ŀ)��(V�����v�oY/[����)�.��M�k('삌�������u�n6s�euQi� 2�>~&�/�)F����+��1�)G�H:nC�գ8Vz�S��j��H������-���>k��ސ�=���R�b.u���*`k�m[0�����D��d��/��*����u���/��J"$�7 ��)!uSc�+(Ү;F-�:MP�>*�����x�>l>s�+���i���$=�̲l���~g�a���T0(�X���+���t�[�h���#���y���غ�@U�)SvX��g���X�cJ�'S�E�v�^ֽW���Fb%�xu��Se����pFq�d�vMH�-H	R��Q���dR�;&[��U)9��*$���$���U�9�����`�=��/U<�y|Q�U���i�p�,g��ֲ�����I�-�d}{/WY�j���c#�2��\>���#�B��"w
M)�L���&�3r7�H"Y�ifZ��c5 3�H�w<�H���YVlr׈�)��WȃR��.,	�ʢ���.J�H�ɁӾ9��t��m-��O$Ny�=��[zd�CWO&�(�ug��E���/~?��:t�e%ʍ���q��dT�,y��_:���� ��ў����jNiL2��Ȥ�9���#����L���"g�,}�a2{�8/6��Ӷ��9�%�~����>$�d�S ��VW�����i�����q�c�é'?���~���s�?�}��s!��+�o���4�ɾ��5K{�[�L�O����&�����vG2�.������U1P�q}��2���}2��U�،֯�A�|N��I X~�������ZTLmܜ}���Z���	@o�%��#wR��=�6+�j����,OR^�i&E��z�W�Xn�%O=�{ʃ�T�q1;R���+��]�u��Bm��J���+�,h�F���)&+��(z��t����Gy��<�^x�_�1�YEMD��bQ�׾���&+��[4"�e������FnJHU]Q`ˑA�iE;�@��2_����Z�'	���r����q�\F��u���
��4?���H�@.+���Tdrsժ�����1%�\�V.	Lt�U˪���r�e�H�����7��ї?K)����&����j����{��V���ūN?/��TL��^a������SY1}��8`�*��_^���s���KP�p��ވG<�^rr��ާ$o�A���;��Ks�5�hV��+߾�=�kؿ
��ه⬏�t?�~���?��{��:si^s+𦷟���̊Ԫj�����1�/��9䠭�����OzN{��h6�
���]�s|���K/�
�Vz���Be�Ń�\�a�T�R��dU�HD�(?���-?H����g�k��2�Z�j���.F���\O�l%A�Pm: L���xH6b�8ZK҂0��̤���Y>"���F2ѝNL�#f *�*;4�1f�k��SfN"�3Z�s�G_�y7�䜘�Z�
�rǯ���a��D��v��詠��,��`������Y��#Kk�!=�,�U��y;�CҤ8���ckd����`���ݻ����9OLӁ���Za�6�Z,�߄2^_�M1�j�A`Z��
͙�D)�C@sUe|c�w tc��K��{4ϊ)�i:(�pK}�4r)��Ō1]�`�ֱY�(J�+��1���g�*� �zL9O�SJ[*�b��y꣜�-��r�$W�5�1e�4I�4/�e�.o��A&���ͽ'�G��5�i��Iy���&[F��́ԬD�pY�q B�?��x�~���l�Qw��8���%,�5-��X�M�"���Q����{w���o��[�v��>A��E&n6�)ʛy����e�	e8�Qۗ�8t�"�.�f*qy��U��)]��"�i������=m���}X��6P�5���GR�v�]+����O��zҔ�.�8`�1�x2W�,��^�מ��[T�}��� �2�BH�$�%7I�����:�ok(\g�j�,I�����H^�ύK�\y�*��C��?�zk��0�N�35g������������8�^���DT� ���\
�AE�3�f��&�4��DP�gI��ΙH��9E&Qr���]h����8���{�Ԝ�f��Y����ϯX��?w>���b\܂��]@��r��B�,�@� ������^�ׇr����A�H�JKFcRT���9�Zu:VG��jq�*���͝�3�@	It    IDATr��}��{����5U��݇�j��h$G���n{?f������x<���˨�]uܳ�R�a��u��O\�/��St��~q�M�Jj��Z��wkѱ�`\W�8[Cu����~�g6��D_i@w�W�w�Go��L���>����i����.��e����h�Oj��� �����"��Z�0U�s�,���Gk���Y*wK��řl���P1SHz܊,�GN���1��UZǟ>�xޓ�-,���Ѭ��~���䍸�`V�
�8����,���־䋛::(k4M�({����8rW]�a��A�ϊ�?�o^t=�han��֖-���7I��X�ؽ27�w��w��D^����L+%�LkU�aI�bŔ�TM��Ru$`�"`��~V��L)/�u+��0�:�Zf��M�>�+(�b�][��}��\y�z5 n�n��H�P�]-�P�0�}�j<�+sMUL��r�*������G���_���k�la��m�6^���2;�N)o S����&�=���+_�,�\��=h~t�ٟ·ϻ��>��7����G��ԁi8Z�JM�)J�pE4�F�?g�1�L�O��s���`�S��>�f���[��w����N��pV�{��}�ٸ�GWcZh(Alր��Uv����Q���c��aoG������������y��L��	Uh��x ����� ��8&R���p�/��1F��OLIS�8���)��0@��ϡ�j�R�Zb�2]J�hr���_�&�Aw��js$*.�0��O*���pj��6"����r�K~�S��U�}+��$V���9�HH߬ʗ��������F(r�v`ژk��8����0�	&�G%fDb�GY��$���� �ʄ$�֠��W���;����f��9��l(֫7�^<��ƅ<�Ȃ���qf<���	I�|�uȐ61�!,x��^��)�M�|?�;��5��|uIy���l�F���$��6Һ��+Ƕj�θ�f��7Qݶ �8��؟���P�[i S�p���
�E���R1I�!��`��i�Lg���`�@�Iy�����f�ć��ds����uGc9��Y�� (�^0���4ʀq+@��:�{^��!Gc��&6�^?m��P E����%��?H Q!HC�a��aw;���?:=� p�O���-"���h��օ�+뎀o�������7/A���*%�i��b�K|mV���.?h	�>�x��[zY ��d�����(��i��{߁�ط|����>���k Ώ�R�Ge����Te���H�|������ȓ��T?�Q�`
� ��&9N�|~��n�4�I��U�`>c�w�� ,E^H�b�l���ȋ�m+$�!)�
Q������q�|���ۜrO��������tJ��}���d6��̳��=P�w�Z7����A��C��}��F�#�*i��I疽��0I��1~���U`���J�y�S����KYsǸwI���� 7�>���7��Ƭ� 0U��Q�Vu>�����r�Y�%�m���=�[hk%*WU����z�V!�a�8p��q?ui֪�g��Es����9��Z��s�"DR�q�@��Z���GX_ُ��^��`���p�{�<��8�`�i��6&�s�Tf��|��pι?C{�¨<�i��	{�K}���*�¨^)��i�]('@���d�9�$�+ۻFdQme�Y�3 �[ ��X�LHcDB��2j��F%_�jӨ�����S�8꡶ dOz��ں'a��� ��� ��e�F�Oӌ}�n �7:����,N���� �L:mgɌ�c
��V�P����4`����s�.�r/|���WW�bV\�tF�³�=��{/��(��z�D&sm��P>�E����v4��Oo����k���cR�N�?��O�[߿�⢀isa�U>���yB(f����]�%��0�2*�y�GcmOV1m��w�xZ���[OP�8�j��*F�6:++t���<#�,����	��~����jM��R��~VLו�+/�z4���L��BA��Ř�b�M7c��rM�#�
0��-Z�D����œ�\�����a{��W��p����Y�?��B��@`ʊ�M����_L[�5<����?~&v�8b6������.s���"�쏞&`j�?����cR��yFӪJ��)B�����y���W`�S��
���M�q���x�s��� �����o�.���
��8l�N~��S��R���M���y�Y���_�+��	s��(�[س<�/�؍u��1Q��_:8�*�ow�c�֏�$�MZ���`&��8�*���5G�*�VI��P;��X�02����@0IX\fj�X���,V����Y�p��y�K��T��d��QL�dv�Zߤo#xf�I��H�EiF$��u`J�=e��vӱ��`�5G-�}v�Z�b��bZ��s�F�'+���'����ذ�!{H��8�%��gb��S���u�`n�n�;%�^M�a�pN>dI��;=Lx�����K�II�WL�2`�Y�b6�Y?�0,��U��
r3�iI�A`
��n�,K��0���y�-2��)���ȥ���@2ι���wQhTL� ������r�qt�*���s&��*[�1v)�Z d bkV���(����1�t$sс���5��j�1U����"=<�#����@)A"%�b4�\Һ�Ң�%J�]e�_�Q��x���bՒgo,%s<��.:���ޏ{�u	�z�Kp�NK�Kn���"�Bk'K}Ǒ��"��v����O~�G8�c_E���=<&���X�Y�"����g=<ꄣ���?��0VU9d���׷�Bg���-��j�x{�O����ž6ӖL���>a|����[P)��B�I��?���	fV�I{U�Ы���J�D��#\�R�TS���7�J>��;�J���Ƌ��ɥH������d奝�����NO�M	n�#K�P�Lz�9�  �%�; ߬7�H�8W�K9�'L���"\�Ӻ҃��i�3'�"\��[C���Zyo��>G�K�{&���&���u�ml�Op�#�?8��ˮ�������K�A�ZϪ��������žN�ڢ�Yp��i�ZDErt3M171&�yn�d'��O�ݫ*U\`�R� �F%�|_)�ɓ�H�3�D)���S'7\�� �?��j�������)l�����Q/�p�#��O}$�����C�hd�����Q�+���ˮj��_�>ν�2���T[�+(��0��)��r7+{�3��f@��I�;Se�H"0E;/�ܹ6��^���'brS"�{*U��Gh��)[/w�YU<{:�k�Z�ŧ�!9�>�'�"�GS�^L9�&�Ɏ�l�9��Uv�P)D&$E��DT(��Ϛ�1Q�s^.偑���8b:�Pb0\�B��W��(<��0�Y��[�x����O/�	(-`4)bDIl�Q>�cÉX�,L���YA�X"��V�1'���‥�r~ƙa��qE�Ə����-&��h,Σޚ�b	�gX����d��&Su�)��a^n�a>�AF�~��X�S�bz����t�jq����a������S�
1��,6�b�]�y3��\�*9p�&��m�)K�4T��YG�LW^��S+F���[D�+����JҸ>�B�5�Q7#�����܄_�M�{Gk�
}��Ul+���?x��i�bzg�X�����X����O| ^���0�����/���~g�~�#��w�V��2��W٦�VI.q����9妶ft;��9����������f�G%tV�1�0��6��;_���ڑzL�����O��Z{L�8���x���ӟv��kv3JL��ٜ��Sܲ�+�F��J��������??u.ֺE�"���Jr<��m�p���^�b�Ղ�_P6��%%���ZC��9�B�;�0�hD�ˤg�j��C�m,�l�]/F�����=�$��k�U9uuM��(�2
(kd�$A��&�`c��$��dc��#�6��L�$cLF2BIH�4�Q�z:Tu����ù�Z����o<b���ֽ����k�-O�`�=QY�9�ɸ���E��3��3W�l�:l	����R�8C�ɒTN�j��D�	�bZ �)d�i��ǴUk���:�����I���d� �Y����Y�%�VI�W3�U�Xt
F;bU=�w�/��Ah�rDɛ ۘ<��]��qS�V��ҧ�����b��Պ�nc5?p`�\���M"%H�+Y,Q"�5��9W�M	�)?V�Vv�w�<A�0���+o�DҀ)�)5�1�LS��u�&Q��AarB���a���d���>hŴ��#���L6��xI�預Q�#3�R�:RI@������H�Ձ�<���ۤ�q2�y��,t쑂��PF��\�6�6:���kJ)SvՁ��c��4�|2���/��r���"�M��XF�:�agg�|>�޿����E(��ϰ�> �I��ʑ��4���~p#>�?� 5��; q����v:��:�Qb�_�S/:�{�UX?Ä�g �G�kהM<��^'���H$A����׼��2& �)�rZ�sƜ�0��Z]�ٻ��P�+HbS�h|s�+��%�1�㮨��͔�� ��#�&��N�	K<��V^E����í��A2lyO�����n�#��^�<�cg�h�6�#�gN������~R�,j�p��Ϫ @��x��]#��֯���|�.�t0�G��Y�S�h��I(�b�Yb)�q����a{��2�������]��N���J����$k[��o�U�_��~��[q�֝h��H�� �K��9�N��-��s��4*7�Qn�j�;xkeƁ��o,����}cc�&����ꎈ�\��l��e�.�r���4%.��zU��֭!ѫaݪ���q���sq��0�Q0�� R��	��׭[���n�o�Zt[͏�÷�8K������(���׊Θ"!�t1i��q���L�ֲWL}�����L�D:l�j���\��D�;�{���hg
i�F��^���ń�~�\&>3Y⊁�?$��5"9��J�z��E�����9�AJnl�T�e�)��1�r�F����8=蓜fKO�v�:^����g��i�3��E�P=`Ǯ
v�]F��P*ok��������|k�T4�g��C�f����Ό���3�1	������#0}�ۿ��nهnj
��q�Ɗ)j��6[��,��E�n'H��6���T?�}dO$d�z~r\�u	�ZT�9.{{8@}Lr��f��Ѫ�b��֥ɉ�rIM�Y�C��7�A��;�6+˲?L��cHxŔf�v}^�.�+�x.'�G���8�ʔ�SU:�����vދ�L���O��X1mV0�Zƛ^t���r�K�Xq�	0e�q�<�~���>���겳�7�z>f�2r�>���鋸����jTq�����}L$��}0�o6ݴ6n\�O���@��Vo������_����`�nR��V}�-0}N�4+���L��O�w�߉�J�N��+^���9c���c�*K6�d�{}T-��@�PD.�d�`�?����/�����I����p+�|Ǝy��@�˩��b�!<�)5�!��HUF��%V(C�"Zý�lH��@�ɇ$NR)�R�_���t+�.{✵6P�L[�`��5��3���l�:ii��e�IВ?�K�X.!�ˠ�jci��N�=&3�S(Z��F=s��D`��*����4��zF�����f�{�US�@� ���L�/A,J ��� S�Z=��Gr_(r,�8�O�ÙW��j��_sQVgި
���!�)���� U�J�&si�2�J��u[iڧ+�?�n�-�|�x`�KHM�O4'#�(#��e�PB�������5�����Y1-NM)0��B伖T�X��A�ธet��sn
� Ɛ�Ƶ�C?��R�.���1�h��bϩS5?ҨD`*j1��>su�����:���4}tK(%[8���X53�U3Sh6:ػw?�����X����I��.՚�=���wͣ;("�Cވ'|��Fr�ը����Do睶��W����㦁1�����0'OdK���2������a��')��ꦞH�Q�����jZի���7�M�}!N�X���	��h�Qt�L��Ѥ�V���^��c�u�3H��'E7@�el�!1Y�H=���?��%-��Sqdo�a���"u���$X�W+��-�6@�*�����]0}ē���98�e�W�ی�(,��zS]���1`j'��K���*��=�Z~y,�=���V��d�1Sx�b�k��+�'�Q|0�ؑ����7��y��L�I0�)��Ry�w0�}��ȓ|��*'�3�	3+Lt�lc���*��
Nݴ�|�8���Q����b� #I�wV�����}���o�O���w,`�����d� �(x��9c<�CV��^�A[ƾ�#���T�(�C�1�d_�l�^5�ϮT�5�/L��V�7��H@F�J��Eᡱ�$�Y�jm$���u4*s�$Z�(����p����	睌�3�D_c���-a)+)-�[��K���}� �q�r�RAMg�r�K\��w6)�f�����I>��\մWח�V�B�[?x��:vPm~�y��N@FnD����$����Y��؋#;L�SH��X�P�����S7���U�9$V�Z4`��$�Ԡ#P¸���B4.�$��9�M�s/�1�!Ib�R��W����3�Ѿ�v{	��.��9������g	[�T�'K�-e����i���X�{��p��c��]���=��9�^󿾄?�~fFf�f�E�A��2�b�Vf]���z���vj%�w�L&�Q��b�NK�D)/�O��	'�4��\��j �,D���S���Sk���L�=�������B��4D�,���@���˸ʉ�`��^4��b�$�t�(-[�D_��E�h������'���'�t[u��6��JV��<W_q���a��Mq�ʶq1�¾���onيr)��R�����*�;�x�G��믿C��6���x'6�s��U��J�~������.O
"��uq]���}���O}�>8�Π�t*/���<�%�t�4>��7�q"�U`��!����g�r�C�TZh7+X�n/y�S��<��I�r-��e�'������퓉M2��?��쏱P� S��eA+�6�N��h���q����o*V1��6�u�gx��`��-���z�1�al���V9�9(�E�JE��4�lGc��8m�	6<�iu{4��y_Q�燁W0���}XqFRZmi�3-{�X�j)ߓr^�4^�,V�mu�gB�����!���}3�p��C57�j�~����kE�Cԗ���@ӞZ,I������ �>Nx��9ṑ�km��3��<M�'��X�b:-MhelNd��ϧ=>:�\�����K(��t;X\���T��]����s� �S ��<2.f�G�U��q�9��0�j�R�T,�C�xMպ ����@yv�S�[�>Ȩ��H5�+�u�����lˌTJy�bZ°�yK0�D_,�TfƏo��ϊi����[���@Lr�ж�I3+.�>Z�E�f/z�Ex�yGbj�3H�NG&���;e����4{��
�?߂��6T�\���$))��ڍz�ŃL/:{#>|�+��0�e$,�z��N�2�HA���R�b5G�5�fx`�!|����~���5��i���f��u&�N���n���aÚ"�q��x��.�TYeQ���R򯿫_�~`/o���*�Te���;��_߶��,҅��19eE=�B
�4�f�Lq��+��*�[z�+������r�j׫�ۀ�eA
L,��^��MZDLem�,J���(��x��^��Jl������u圱;�g�V]c�=_1)\�m[��oy�3��<m���z�4��E�5 �SNf(���<j��Ty� F�}]D��5FxvB&����5X�U�]#݆t�e�[��~�f�x�S7�K7�؍eQ'H>c����
P�}`��������c_�D��ق$�|$�sH}�    IDAT��f�-'J`�������o�Uy�f}jp��Kã|A[.��q��p���M1��$���r�v[�͖�k�����A���8��Mx�%gコ��̤���J�iM�%!�j��� [��{?���e+�U�N��D��T�s��Ny�xeG̃I���j�ڻ�y�zV�2��N�<�{�G��cUܔK�'�����x��ۓ�Pd��xf(�X��Ǉ�z4�3�׺�	3�#�&�U�l�c*��Z-�4����%������y�""��qs:����3D���P��ZbF4�����{"���q������<��^����ٞ���dd��.~gյF���L���V��l�~�߷�av�R�\}�^R]?���$��� �6���佉���DO�a�51;>�d>��L/�zL�]�$~S�&L��X1m4�nu��4��	1?R)�:��"�2�A,0��P��G��\/Tr�b[*�ҍ�D�!�E�U�R&�q�o�qh�n�j�� L�ʫ
7����6�Zf��E�֣#����LT񖫟������2�>j��[	L������S�;��������756��z
^���a��}�
��v",r��>!e��yN�=H`���7�o��Ժ91J�rX^\@��j¼�k�(R^�1}� ]y?��oކj��vc	�����_����Jl���`__�ޓg}�Zi�^j�� 0@Ͽ5~z݃x��~��j
�\Q��t!�H�#��К����E�"��*��Y��|����a܎V=qsW\��Wԕ/&�Ow��DY�6q��9�z����b܁�/&9�BJ�b��zeU ��۱U(�+N@��G�<&�pz��s$N2%lnu�cF(϶*��^�ҥm�;J.5�j�V5��� �"{/��,�,A;d$P�H��Tf�cM�S3��!0T�`��g��L�������mk:JDe�� m%�S�	�~b��Z������X����Iq�-���hi��f�	��pt�����#��5��à�q1dzǊ���Rʛ@�K��AC
�5����Au|�j�MO�Tt> ^���C�1���2ڍ�>*	�%�'K@�R
,āTL�c:T)/i�z[$�b~d=�L��ϔ���ey�遬DRB7�|��^� �z�f���cͤ�X��:�˧h��V9��~
xx��/����}�Ǒ)��Ya[�
��D�3�������{_�Y�A����*����Z��ZLg�T)#n��:&&�3K3�<2�,R���-�����R��8ʓSR%&B�b0 � �J`f����9���(�R8l��SO8
G�_�r��b>��k���0^.J�!���� �m{X����1�p�Z�
�������]_��oڍ~v���(���&M9�$���]XI��ʬ�k�!q��@7M�������j�uc$}1����[�U���6I��Bw�%,Q,u���j��TWy�Nz�,.�5*	h�h$	ץ�3��ű��C�DsC����z��l3)�WbMu����O3�}��JC�A�(aP�{�.�#Rh;�$. U���V�BOB*�g����z=��l���D��~k	94p�	��+/����Wc$'�c����[�v�d��~}�]���{q���Ic�qْ̓��)
Edi�ıH�K���u�
�g �9���!�h�^��г؋�2j�̼�i�Z�,�IeF�Ԑ�����2U��&}���G����3��7��3N=kWk'���=M��m4��������~���}�"�kC��Kh�A��ޤ��S�$�<V����>=��f`rq����A��~P�ɑf+�	#`�Y����V<��h�HxɃV�!5Z���g/�c~����gMN�j�Y���ր!ٳ&�wG�^����:ѫ���8�P��{�yhl��
�#}UB�A�}_���U���#tR�z�*fK����x�S�	��+;��ʢ�s'��VO��B?	��i�h��m��y�Uo���l"]<�1�����\��T8�x��|�@-5���{���-G�P��9� �$���E��i|P)/�z��9�g3R1%�i7��sT���t�N������u��W���5��Bfg�l+��)���Yq �b����\]y�؃v��=����J�.�=��&.���Xy�u2F�������!0}�՗��gj�T�3#)W�ӑ��;��~{�}(2x�3�`:[JK ھg�k?�%\��wc�O`,�ñGM㵯�
�^t

�F���4�3 j�5ieo>::�v��[�ßޏO|���3�G/Y���*I@�
Z�CLOޤ���cL�b�m��?㦛�G�F6���k�x鋟�?��X;�`B���jU��Q��| �-[��~;�w�΍�41�T!��2�<5��%�l�6��mp���`�L)�6�UD�'B��ףZ�^���k��?ݼȃ��mi�D�	��/�B(��"H��0��o�rx��5i�͋U{��/�޶4r�JBײ^G�X�f7;�IπZ V�|!�`p!	mc�\�r�
�l�2Ւ駶��}m�ݐDSu`֍��X����?��}�j���(�����&y&��26N�^K�d�����`(a��0`���G���$~R5M�T.�Sʳ��i��y�td���Q�	�4g�(�=��h�s���VL�2.�I��a�lT���R^Z��(�&d\��b�F�+IWLӔ������
LY1�Ӯ�,$X(���@���N��a���rIa�l8�TI��'H� ��Y�x`�[Ȥ��k8~Co{Ëq���c�|�dA���^"��.�������>-��7_�^r&���2v#ٝ�e�����K1�c/����[����%���X�f�8xS��s��q�]��{Q��u"-��XC"��b������H�a��!�+h�XL���{�>�9�T!��b߾�X\<�b���C�q-���\\x��X5;�\��u�dE������ā�8b�*��9O�����~��M������;�I� �y�ce�R�*������Q�Bъ��X%�D���&�RP��ԡFB�)&���8PD�A�����g��gq8�!���`�.nL#�[�L�L&l�ԫbTB���I��쌍ѯS��}�~}u1�
cD{2/a^�*~��󅷶��սl��r�c�k����2r=D�z.�,s7lY�x2isp�;�/4��8�Ě����>˒ ��kd�>�,b�LW<�l<�)��k�������VD6K�$+!C`�<�g��~���|7�>�s�6��M���g/{�$��Ng��d%�W�J n.�|1$U#%>oM>8hsG�K{�Z���o$��'����i��騹Mi�M��1h�X��r'�r�)8���p�aՔJv�`�u�+��-,ր�8���w���Gp`��p48�9{��B*1F
K�K�Hz���%��_��(M�~jF

�~�Fg��"]t�S�Tαx�v�U��"�>p��<�ĉ����˹�)F�zLҽ��B���y�q�_�<�9�җ�����a��I���c�m �sǌ���W���y��?���pg��\�>�3&Ryd�l	���}ڙ���O�tV���ԤR�"�%wЈ�ǒ���{��^�J`������,�������`�\��5�X�g�'I1#��G�y�:�X�1z�8?7����u�e{bN*�y)ťB����C�R	�VRJۭ-��0�� �.�RH��a������Sr�%�I�7��mP��e��	�H��I!���Sr�˼{0��b^���;����	s��2�Q7I;b�F�z�͏�0��^�:�EL'�x�K.���R`��i+�X]�aH`G)/瘎��a������k>����{���O��Tq�G����s�Fq��7�T��;�h�Q��<h�@I����x����v/#]�� �E�\�E@���~��<n�>��7⤣g��3v��!�qͧp�-��l��vp�ч�/�S\y�f�<p3�kpv���L&�����H���b�#dr��^�L� �x]�V5��g�����B���ܰƓ���Jh��A�o2MDt�G�{����VV�:1�y�~Ti�+�*�V����7^�T�Y|����R����V���H�|���:��: �f���\���P���w�ٕN�����%3L��ܓ���{8�C���O�u����/��ކ��272r *��9�
�%��\u���et�UH�ʪv����3
�o(�E#�dm�׌js���#��U���\g���5"����T��H���*�L C`:L���`���(��{ؠ/��&S�SJ��3�d�X1�0��e�{L�4j��$��S�[��)e��t*U�1e�O��i�1� 0��0q����/���&�m����ňr �P�g�����O����$��UQ�4�ګ/�UO��橇�1V�V��'kOcH���p��ѯ�{�)�Fq�,�)}��w~n2�E<�	�������PX_�<�}���s�F��Q��f�mݎ������e��ELNM���b���}�v,V��,�������IUA����tO���c���X��;�܅-wm����X�*\���񸓎�T����*42�6��#|��?�#;���u��^x��$������|?�Ճh����ˏ��H`*XK�f\��q�E�Q1��x7�%<ܗtSW���+��"#$U<v�sD4�y���P��%��$zj�s-W������&�~�RZ_�
��g3@�#:��I����[���dzf�i|�΍p�ń� Fd�'�3L�Nqi���:{�'��߿;"�Ԙ���W����S����L�8�l&m�����Nʰ���7a�|�	�&��:�C���x����+����$�P$.ZUL+��GpJ�H
hu��
s�9���7᷷nžC-t��e$�C�]�sP$,RA��)�M#+�Q�|MF#��r�WX���F���گ,�3^����.�������!=򫧊8� �EO8��-�(�K�o�=���5�a�ۜ���;?�?��;��Pm�O��Od��k1�x:+�S�29X�7	D^'�>u����|�'޾�Gᘭ@�1�`����\�r��M҂�w�)�-7T��#��+��D�_�!�Wpt�A�"w���`Zc��ժrP��9@X��8Xw2��33G���[^܉o#u���"Y�����`ᤉH�U�b[̰�b�����y1N9zeM���л3���Z�9���u ����Y���Sdk܆�H}`_��_>�/|㿰P��Ƭ��$L����v�J��!�S~o���f=��&�b�\r*�M��mPg�Z>˖�$D�;�>NJy�u\+���NN#%�Py9���Q�p3*��ʛ`ڜ_���H��'Q.ɟNJ{^]�!fM��(dҘ`Ŵ���.ӦT[��"�t.�#����x��G�|�nG��}�eO-�-/y2^��s��hT =�]�ao�A
���z�'q���G!�����|������}>�x����� ��!
yι�"�
�{��x�+_�SO���J���c�0cVI��,�2����_���@"7#27����1��U�Ь���z�,>v�p�Q�L	l������	�t�V�j��I\p�I��W>��E����qKW���~(�`��ϼ}W���Oᾇ��HP����H�h	Ko�4l	��I�ϏA�����S\< I��tu�xҠ�p��=~P��V����zY����"�R٫��hޤ���Fc�Db�	����p	�-��̵�7C�
L��b�gq�(`�,2��:�8v:��;@�ӓ�={%�2�h����BR�y�W�c���t��#�-U�V��ʌ���bR��F[$�V�	3ϴ'�ݒ�^k�V�9�e�i��؎Fs��@KRM��`̄K��H��)�k�!W]���A_Z��^c��IjR٫����S'>\��*"�i�m|L�����)S~����'CY_e����S`ʽ4�D�sL��>��{.O�#ѝ��Z�)�iz��~!���YodAQ+�	��R�+���@����U�u���t�dP埢.�
���+*I�﷿�Ur�j����ӓS8樣P�,w8ġ�E4�-�^�F�|�*�]>���{?���Z�O�ꘓ�Y��w�C�����w�S��ZR�]�h�V�KuBD�l����u��3ӫ���gEui��Z����*��������"��٠�\&��f�jf�^K�vw �����S7��q��!$����o�'��[�Q���_u1�Lf�3��J`��k����b;:LeNZ&kΈZє�2�,i�����"���V����讏��:��~u�U�/2U=3��#��5�'��Q�I��<j�vsOL��:f�>Uo�m,���NB�!Dw"���O����=���^OB�'s���~��獪9+ϊ���R�*L�U�h6)�$�-W�!1���I\M�ݡ6J��_^�kQ#�c��g��6*�cZ�w�/��R=�����G���A��Z�����̧<z�y8��u���F�Q�A5�`�N�O�� n���|����.�ۻ���C���j⨪��qn��6��ۉ]*bTb���5�31�w���A��F��@��D"���X��cX�n��Z�6m����7�09&ܠ�����h>���W0���
p��=���o�o~��mʗ)S,b��"�f���ִG��pL���	Ezo�+'�t�%7>�Hc��#���<�>c��4����I� ѕa��7C<��[]�J2Eq9����Wĩ�G�?L��+Ѿ��3�cQ���<�����1��T̊B��)��6b��hk��*I4B$�d-@9���5���맋�)�1=^B.�B>��sF>���(����(���y��M���� ՔtlH�&	�*������b�B��e+�[��\aYq�7u�I˵�5G1�w���iV�����޻`��K�x�`�)M�"0uO��X1M��|����j*0�֥�)$K%�񊫶 ��b<3)��B�Т���!^T�qf|����c6�HȆ� SVm�ʻH`�hI59[bŴ�>e����|�1��������]�r�A��~}3i�'��:W*�LGw����UL!0�����m(�xޟ��׽⹘.ho�v���v;6e�G&=@�1�B���6��S�x�r�9�tĤ���(���c�mp�,Ə��w~t=�̷�E�ɒi�H�fP#0�W"ٯ��f��k^����
�����߾�p����jq�P��9ox�qṛP�`���`w�� �\B��)�X����1�x�X7[�J`�� ��7~[�B2]��[&0L{�����$�I�(�ݐA��=x
2��:6�(��X�p���wEJ!g] c���>R �5��*�D�`.n�Jh�&v�<[��]��yrF��&wQ���NH"e]$�aSv1�l.�3[y�S��n����J��0� �y[�o"��vM#|����!�MK�l�0eM���k���+*ya	�����h��@��C��ɺp��;jɗK�FlF�Ci�\%��t~��Ԁ,��3A�o����3D*�R����R��^��.K�(g�����V%}_�y��صx/���V=\*��&.�LHŴ�������#ʾ��i����)���]���L?9��:��&z�e��m����1��)a�X�u���?���H>e3���N��4���=r0eŔ�^	VS��$��6�q��q\������گ�{���A|�ӟ��M�pՕWb��?�w߃;v�IO�e:�P���[����[?���jL6+St�;���<�v�q��5�ɬ� F|��h��F~�x�݅�7��}Ş�v[J	yﺜ�ʙ�29!�~Ѡ�����lF��5]�Kl�x8�<b} G!��#0}x�?¾K8z�j���a���T8��v�W��_=�vr
�R��	q�n1��y��ZY�^Q�
��j��ߘ�h��qp����N�p���؈��EU�80�긑C�|ZQ1��:�fF?ky��˕=l*-v�׮H⁑SV1�{�6Y��B�j�[��*    IDAT��f��J=?TU�_u��g�����*�`���JM��z�7�PnƖ�\.SՅ�W�'/���y;� Њ6j��h$�qi������{(��\x��y��z�*:�E��ul\[�S/:�x�f�p��$���=�^�Wn�{P��Y�i��m,��m;q��=��nl`/���hS�ec&��!AF���`2���3oY�0?��J	>A�L�p�q�t�t�{8���'��Mkq�q�v�8&�U��Ń FVH(���x.����t���߄�n�{��E�TIzI�e��r���Ǽ.�U�E��!�*��?���s4z�ͯ#��2鹥OV�Rݏ�C{!�;��N}?��^�������qIr�{3�I�O#�ɣ�(���!WL�� k��j�t1ɲ�4����.���X��Z1��	}�\ï�`q���T���Ѓ.g�����Eu�opQ�^[�O�u�w8q�z�c�ol�y!��� �+�^�{"��F�����,�������,z��2�"�t��d��2cQ�,���[�pC�Kh+u{4���3��dެ��)��9�4�A2)�@��#�=�ICdC���TL�K�"�m��P�?>)�G=��r$���	����͊i��y�=�Kh.-˥�b��'��.f��!?g�{�tPoȸ�v��VV�m�����̜)��f�*�����5�"�A}�ٺTL�cʊ)%��4�)���H�}}��?��M̏L_��0[LKB�� ��*���AT4�ɡT.P�Ak��9L�8�58儣pΙ��������������=s���q�=�۷�Pm�Li�aY1�:�2x˕E�1O��p걳��5������ج�r>�[��O����h�"�o��ӎ�[_�\\�''#�j�>�����K��m:��F�-�Dhޱ~�Z��˞��.>c����o>���އt���U��#u�1+y�^wv�~��\l+���7i2��+�H����z#GO\{��J߁'s�;�nj��\V��� ��CB�x�k)��~	a��K>�T	i���"I 1���"�f���p8�:R�LPJ�}�nd=6Ы&�A$ō�m��� ���W{���ɣ �=x��d����遱����)��r(�<5t�C�ׯ!�:Z�tC� s ��э�g�2�"�
=���.B净��FٷP�.0v�"ge0Ns�搰T� ���j�4�i��N��f�i����S���s`�aqq	CJ��\L��*0[/�<�')�7ѥ�O�-.tL�71,�ѣ<�eӞ�0Y�q����BŔ��@L�k���<�Cv0$0�<�ӏ��{��<wxF@/πN�Gw씵�n�乖T��7���F&͙�C98.�ڏ~���;�)�Eyz���*s�?�ˀ���5��T>s��5�k��hTj-<��!�LL��q�J��m7��e<�3�����͒�w��Z�����ON�#_��B������Ai�q�k?�@̓C^��CZ1%0=f�ax�b�4+�L��ko}�W���E;�R^��3��cI�VHm�0So�0줊U��\7��k2���+ � ���
z-����niel�垖��y����X�}*����+8�!�n��.@+�����T�X���aOܼuƒs�O�ko��:�?��^籑g�_�~h̐6���>YǓm�W0ɜ$u��mH��^ �P3�b�2r׫��ZV1�:�5t��v�ɭ�"{�҂�.�$��a|�AG�a�%��IHS�~��^t6?,#�J���<KZ�������:�Z���G`�#�u�C��v��/��\G��9q�7C6o9P����=$��t�\���<���ذ~�:j�|�	8��T��ӄ�6��b������$ ��n�?��ly`?*-6�̲_��ݔ���Y͒3��_uF7�T�_=�d�X�I��;����x �+��V�E�/\����[R�8-LZ]�/7��~;ͥ<�\���H��#\s ��������� �^^� 1鹍��;�复�4���җ��R�h&�g�M�� [�(G�N4�A��r��F��n�6���	�r�6���h7k�q��(
]���oAt�'iA�����[�E�ͥ��}�`I��K�,gd�4��n*Wx*1�bȢ����M��;S-����%m����S殁P0�P�����q1���q��z���Iqt
e��ȕ��GL�9$�'Tʛъ��'!���'F*�2(f	L�hZ����9s9d'�Nˋ@�K��m�-�[�R�&�y�ڽ[Z������)�y<�S��h�J���@s9�u���s�]Īlo~ɥx�g����|�'p��0F`z�VL��:��}�{>�5�p�CX�����<�!u���0��av�/�X�H��X�kwzh��h�B��B�Þ1Z���H�L�t6��H�T�Ȟ1j�9.F��>~��q�QS�o��wOoz��[���Tg=���U�Ɠ�p��[���K_����Oaq��6K�b��]w������W>Y�)�!�����/���}H�K�\���<i*�$ș9e�%�F7N4�D���<ZQ���6�&��>+�]�?k�p.�P�	�,�986&\\lS1'_�l~Mv:V3��c_�W���1�JR����r3I�D��s�<2�EI�?�k ����RJA{d���@��\C?Y�M�mL�'���g�oՉ���{�R=+�l��I CV�l�G 	 +�(N�`?��Ú�\&m͛#皲qݙ�pN�ؒ0�RzLU�&��C�,IŴ �Z��Q�c@9'������R�T&P�u����۔�L�#=5��)���g}(:~�c�n=�����0���i�1-��H����j=�	�ڤ �A���BE*�P�$'ƥ��KI�?��^F!Z��+o��ð�ĐҔ�Jy��G�"�JkVO�!�4.���ZĆ�4���?��g�1�ӛĚ�%�X�:����MD�4��y�����A�&7h�`gRX�?���~�sO}±���^���(0����T��	l��~�ܹ�y&r${��	�r]dU6O"��Qγ������
g�R.<>=%�EyO���¯~�KLNN��/�Q7^������Q+�_��a߁
�Z;��>�Bl��J����u���e�솝�g�-��0>��$�+&9�����u�`�\y�Ьߋb��z/ȠG�T�<t{h�v4NF���9��cc,FL�,�՘���U�L�O�&;�%)q�ªj�%�x+��,GLk�p�GN���σG��$��/�Ө�j�U�L*M��X���N��'��+�p/
�Ne3�{ڸ��-����1���a�qy��d��Y������~h��W��2�Lho9�n��{u�[G���\��c6��ٗ_��/x<���Q�Ԟ������:��\!�O��~�ܚM�Z�Zk��RsKX��[���V�3p��M���CS�Kx�DIn	����R�tn���X�U�q�iq���K���>q�ܱu'��W7c���b��Y�q��0�a��{�&PU�s�9��.*���Qr'vFF��P`F*�J�V��u�/�[ysf��ܼ�6�I�*y�;��[eN�R_��+#"V�U���K�£3�*���*ʫ"�����2U��%�<֯��6��=�r�򌭥!V����ץL[��)Y�I������}A`��$\���ߜ�.�D�'��qu=T��R	GO��x8������gЧ$�ơH�[
8$��u���Y�I�#"��5��|o�e$oKp$$+�������Lj�汚�C9L�3�%N5id
��2�/�� �̕(�+/{L;�զzJf	�k��JŴ���Z�{H�3W�q1�$h>��>%-a�4��t�gŴi�|�q��J�T
J䚅�80m�஝R1Mg�ȗ��K��K�#3v�ʰ��&}6`J`O`�vȸ�򾙮�L9m�1���U0?�WKzLw׃���W��W��*L��p�������q㭏`a�'ͰS�V	��̚<�^=�68wrY�:M��md�k���#W��zQ��H��2��	:g!�̌A0�}yP���~ܬ ����������o� n�i�HdX�=���^�8���m�7��_������s���`z�1G�_��h�i ���ϊ���9�n�^$��Xu�8T��:$��W��Бi��~"�=^�VZ��rp! ��-�s��,)�v�a�X�1.�\c?���Q*JV�~0I נ��4�o�[�K�<�I\u62�5�U��s%8���9��OW湩|P�uɬD��M��@�J�3�����Tc��p ȡ�w�A�c��<�s�S�yc(�L��r����Z"�?뇀�/	�T�ևV!.v�Q?N��}��y�ҼD˘��a�)�0p��KLX��D��C��ԍ�D�k��nO��ns�o��(#=UF��Q�bQo�n8�&G&��C{����!�m��S(Е���vI܄	Ԅ����4�٨�1]�bHy7���	L'J��ɓ��UA�ǝ H�>��.����g�2�TE$�f| ��L���ۭ#�6���{�s�i}Z]y���<4�:}�T>��hW����<>���㡝ud��HIu3'ӥ�X��+�����'��Z�1�#�4����f��[oۂ���p���7'�;�>:�T���d���T�ѐ�V8�_^C�k,��X}�����c�˵e���{����f��1h2
L��;?��}����<�����}�}ľ����췻�MN�P��ą��	�3{���U��� ��w(�n0#�>����K�ul���@�������|��".��/ֈE�^�Y�mz�W?����P�~���-^����\�h-�/y�/��ѥ��+�x��d��#U!hV�L���Řz	��1`������<�jzOI�j��`�Ĩ�6���!��R��&Mϣ��I���2��c�Kq�����b#-Dۖ�i�Ow�et�Ƞ����3.����p�1�0QTp��[_����_��K����AΌ}���Ð��y��|�{:�v�~w���rb\���6e�y�18-`��~�6��-w���w�`��Dn���Y�9�5��i
�����~�	%���}�����.U'y3|����d��� WN
Pe2Q?����<SݸGe�&���rrNűN������Y��_�'W_i�8 �p~9���%��F~e������]�|�gm��{��?��Կ�������@TRF��s��%鲯W��q��O�	���O�d�h<f�3�t�f��-�aeO�lm�Y��P�=l���g��4�k�Wu���=IM*���x^���fsʝ���>)X��F��4NDpI��'
"3�����`ʍ�����VL��9�q1S�1m��?=1��X��g5��G1�J/.�i��V�CR1�&0��7e���jqMOM�v)�Ә,d
��ΝBR��L��t�$-��l�5�Qv^��`,��,�&�Φkx�K�,�1�1����3�X-�{���;�߁�X����_��lF$�
0�n��Q���qLLOJt�VG�Đ��1g�����ʪ�2)GH6ɓ��DX�t���z.TƘ	��P�}r���%�q�a����ƀ�2��"���ZCp|�i'm���ꙸ��Q�a�@����С,U*����xMMM��c��Ԙ�����~�U�Y�v�~dK���En�����2s�a�R��E%�l��m���eZvO�"Y\Lva:ng��T�!�Q~�@�Ԑ��Cٞ!Ҕ���9�꺻�T`�g�|s�u m�_.Ӓ�R	Iye�Z�P�mMu�M^��K� G����~��v��sB{��h�=`�cٓx�R�'3�������`O
�>Yb㔯�)H����2��'U@�H��n���:�iF=�$��P���֫8A�(�1x}�4���SM��c(����XYZF�^��%6Z9U�K�lΕ,+m�*&V1%0MJ �!�}���D9�N��E�*U$z~YdH&�ʛ�����0�Gi��3�\�&:KUZ��9D�`jr���8w�\`���)7٧ʊ��5���e<մ�rg�S4A��,�')�(�� �N��.9�qx�Oĩ��`,�����u�fTڣU���_�O��w"��A�4%�P�����A,�t�p�G�x�c��+�s�f��n�
�<�9�t12�d4��c���`�'���K� ,��k&�Hw�X [���ԳΔ�e�a�ʡ�l���oǿ|��x�k_�s6_�@.&�i'x����{��h^���X7E`�ʖ}u�1�~�۝LK��2�T�^��y'��˭I���U稼	��+R�Q$��Y���=v�Y$�(k���Dct��	M����^'�Ӑc����N���0�c��HԌm]���j�v�Z,����xu���z�� �A�ʀ�L�T{����-	yl���q�'�l=�cK�[��=R����I��$�se�2`����
��
a��ǚ��}6 KS<h�;��H[�>Y;�#t�6�3��+Dk���A�����e?\�SG���$G���8q��8��cp�y���'���1ͱg%��H�Ý���:y�zv�D���X���B�'ۏ����n}�47�̡�~��'���Y�]lt/����=���:�J��z7�^��V^z����G�Rx6��B+���+�~�^Y�����j�Aw�v���*�4�O���\��2S�*Y`��Ю>	rMrV[��b�+�BϲU =���f#9�G���c/�-G;�#"9<�уݫ�Z��j�����M��� [+V1��rC�P6Ю�΀�H﹑�n�ϱ�i��C���0��C�jv793#�+v9NN�%�tN�#9�.�W�W�m��|�&��v(��܌�1�<V��z��N��޻ey�����B����)�b*�Ǚ
��B���S��I����Q����Hk yǳYt��Q'0��
�͘/��׀�����ϤR"�͒�����y��	L�Hs\M!�+ג�k��9`��R&��B�zw�F�ْ���R�� �n�/����=f����/�x��}�	t �i��7���1%0U�����A�{w?\ǻ?�)�~ߣ/g�b����j��Jy?�u�|�,V�(MMbf�a���[h�4H�EIP�u%.�gD�#M��+ԃ�����rX3����*��Emi��"RL?�W��#&����l�������mw�D�K#�!69�W��2\�30�⬁(*����q9ֺ��	`�N�5o��l�G�4�BY�(Obt�(�+��׋��3��Zs��S6�T��W�zs� �R�x�N��!O]=pyӾUi� Ո��t%R�㯼��Ec�e����IIpY��qZ�"f �J �Z���hh�Mۥ�=��PlSgRN��J��f��J�c��h�pꇑ������ <㠔�T�p��a��Q���=0#	�:R�9��&��ٞ�i�hퟡʢ�%${��I��8[�=Z�^�E*M4�1���)�*��
0��Q�TEʫ��'Zz%�Rmt�oV0�g�:�w(�m���OO!33.���ƽ����K(Mv`���N�����"56������"w���~�3ڨ0m��XA�Ƀm &�I���R2+�T͏Ԫ��̃B��H�������H!T�,aՙ�ZY�Ϭ`h�V�v1�,�]=�j8�#��_�N?R*�ΗK�.V�}h���&����[?���bq��:|s�,�|��a�TL?��7b���K8�Ö9c3����]�'��I�{�*���y� ��n��˶~E��gĊ��#���v�Z�љ��G����>ͥ�]<�m�y��qꩧ�o��V��ʺ��O`��<���
{�.��u3L�"+���.�b�%��Ɲ�$�P��D�R^��D��0uűTL�ҭ�2.�	��u��<I�/���B�T~����4YS"NM��+R�迈Bƀ�S�_�dL�E��i�:*�b�f�&n+���    IDATV�Fk���5I\	fdQ,�ಞ�B�I�^��s��X"e�Ab��1`�g�~z�D��u���*�N��$׌��z5�	M��%w�G��E�UC�^Űז�G"U@�^JG�H�t���7	�����W�a����l �!_7���3rG��n�4��S$ɶ�))Z��e�ߩaЩ#�6�.&r	��*ᘍkp�Y����N�̤x��Oh��aQ5ұg�+��G�x�W��s��
��4A�K.B��(e�}`~	R����G�b��2jJK2��<z	�i��+)I���+R� }���H����x��I��1�(��=S�_V�d��|E���rUZ�Y�`�p�Q�.�i)p���l\��xK��`��Q�����3i%*ZN�Lt�\4NJI%�!b�%���QZb�&���i5#��KDm[�=�,+d#�7�|�;�g4u��1�����X1�]B!\s�c���X>��P4��jh5��1���~�Z��4G&�|��i�>�'I�v�%�G�=�M捶��7II�7zڢ&����î�hl��=+�8�����ř��A��L��qR�O�7_�֒ 㚬��5?JKŔ��X�>j��g�ĝ�@+�9��VAW^��*0�Iy��'�`�[C!׊�,�k�n�qhJy9��}��1��� mO44u��^�lS�"��u���->/�W�1M�u�̏$��vf2G!��x���'�R1�Lo����Ȏ�?ƫpuw��!��ۗ� @翞}[؍�X/��|���gc��Ĕ����C_�ͷ?�J}���$&gg5PqC�!I�B
I��-�2Q1���s%��V�tde�wm�)&E�6K��*H�q։���w�
�Ł�!�u���w�F�K��#֍���y����X5�N
Ъ|.���[��j���y������]�L��1d<$��q ��>�Ǵ8lv	�tD�k�p���ֲ��Z�p��K��St��jҡD�q��T�aєd���k�}��A췣4&�@�)���X���<�7�~�� L��AHZz�8����}(���=I�(��vH-h0V-��Er�� �j�c�m�����8I�B���5Jc�D��i�7Y�W;�4_������nO=b�Ϲu�3*e�h�h�m��o�=F�U�x.����Y1-	�\�Aє{���:��\*{.����8.f 6;9���VLY-�?d%�y�2A`Kc����"z�̊h?>��Y<*24�ug�?m�����zSz&80�z�|��2��;�ge.�X�7�
4�y�G	���cJ������db�'��P�k�MM��'@���n�(�YDzXÆ�rx�3/�e=^��ݽ��~s+ڹ�j'l:�^|�=z��&��Y����;�r_H� �-#_do}
E��&��8���;0l�Ǔ�;
��țLň'd:J.-Tj��n��'����<\&��`�u� vn�.�I�)����b�f�Gd�[�.*��8.�q�Sqgo	�v�V��]�R�_�
V�Yg�.��-��0e��ȵ3x�37c=����<�Į
�7��<��e/:�I�'Q��2GӁ0܆u�i�9�?)��p�
{]J�_%�Q���36.&ֆ�W��	�S}��̙�*����pC�C��2V=�G$����c���Z=�^��a�$=��ɀ��q��}�_�����Nn��b}�ylt�WfcɟR��C�
����F2zU�$ů����V��t�2�HZ(�.�0^H�����|C�,�	�4Z�B2���n���Y�Z �W<X����J*�p�Q?��m-����DۍP����g���1�td^zr���A��v}�5�nvg�q6�w*�ߴQ�cL�hR�3Q9�Ţ}P�=k0vnD$I�i"�`⹋�ZF�9�z���R�����u�����x��=X����%���ʖ�Ge0Lf��J�4Drc=�JDI^`3I����Uo5b���RbW�H/�Ϗ�U�d�8��0�g�$���Q��^��V]�Ť�-�Q9�QR7Q��#�y��e�f.���6z�^e�����J[��
�Q�X�W?�WZ鮷�j����G2�(�pS�QӦx;RDٛ���qb;���u��\+�?�o#��rS/���{����Q��zud�M��L���eٟ�A����� �!tyi��:�1>K��nO�_��*������� ɀ)ז����R�&����� c�Λ�ʭ��!��ԏ,򹜒�ދ��(ڙ���ZhP��yύ	�Dʫ* M��`�)+�E��M�d�S�����6�~_zLǳ����wEʛC�=��"i�u��=�R��"���a��ڜJy����tC�XS]��"�GW^Jy��y���A�I`��9�
l3�K ��/Z���kՔρjYt�@c	��u����g������ Lo߶��|��q����������W_9L�����;Ee����)L�Z%�$��㔹9R�P�Qec$�i
)D<A������'�M疤P���}�UA����O^+��؍�R1eBt�!�y�?c˽����i71^6�u.{�8��̌P����Z`
��C��E���b���K-����]�;YdK"=f�S�eCم�V��6e;S�.�B�ꜜȼ��}���uJQ�`�z�o֨Z=Ipb��V��V{~��q��JǴꦯ����;dL>.�9��Nk���2~��8��.�|�L�q�^R�[����m��r?Cp�By ��O��tc.�qP�b�d.��J�J�Br��;݉ۢI��ms/��+�΍�4���K���U�*�@l�:C2O��>��u���t6��v�P��l�L5��2J�"���.-�Uoۨ	�EI�L�kl��v���	L�R�&���iJ@�~#=��#�a�}��֡
�t�#���].�L`Jq��5�ˢʌ2d�ėh/TЮ5Ĺ7Y�!EG`�+����K��3�B�R^K��A�)��>^�e�lErEG�0�rݩܗ)9�Xzv�HۨWbÚ���sp������ݦ�_m����C��w �� 'nڈ�|���N�b�\m��}�:|�Gw`��C>;!fD�\ű�TE��xh/z�=��#��z+fK��T��kCCɮ={q�ͷ������zV�dL�"v޿)�0�ѓˀ8�K�u*#�u��D���)��N��2���>n��F|���{���'?�Y�u�9!�16<� |�0�#����hH�$v-ox��p�ͻ���3�����AL����&��R��s�G۸���89��V+�ҽ#n�Q��J��iD.����1���2E۵�9G����A���E*�X`"#��x5��}&!�͵����A��ip׎�oz�W����������D���]13���#Fƅ�5C)�)gH�{��M�*B$�H��.$��)g㢳O��)ŭw޵?��v��·��P^�V?��=��Pȳ��Pn�:hF�vO�FI����INj�!S���s��3P#�1�~G������-L�a�a��613Y�����7��1G�űG���5�2�E)n+L[�7T;�p�\O��˟�c��^�s���v�Î�{�Ў=ؽ�����=�b89L�>�͗9OB�O�7�,A�j�N$�l��,�{��ba+䉴c��ǡ�K�}i�'��c#)�hC�J�i�����5O�e6t�Au�~�&r8j��`�tع����1d�c�'�X���(�X�kTy|,\��#��1��|C��="7�
�H�Y�4�o��+a�\���xN�׋&*D�c��b0��h�X���
o�E��Oz�8�9����dP�y��'m>M�E�\Z�����w~��;�d�,g������1BI����/E飽�r�d��#�z�|�����ͧ���g��&����P7�� ���.t1[-���VU��-����F]zAG�M,��7x}^�Bxc��ζ.�uE���~�~O�i9�A�VCu~Q��̧h����D���L���>�]�6ƤB>�R.#=���E4�c����Q`�?�x �J�+/{L�؍^�+=�T�TG��Y%p�BU���y�t0m ٪`&���~�q��Η9�����m�[���ڏ~�>r �c9<����<��D�������۲�Z�)LͮR��@��جk4lA�H��_���{B0}����0�1��f������9.b���;�p|��^�c7�e!�޶eG�z��q��y�;t�M���0^��f&J2�6ǆ�<���k��f���J��.��@;M�`B�Y�TZ\X5U��%Rj�Mn@�팊�1��\nh��?���dIfENw
���	@L���%����
HE�sWc�M�k�9��0�@���RQ����h���T6-�x�4w��2��zt�m��R�.A)��J;<0(�����(9:[O��P�ʎ#v_����3������*�JR��+"	���R	�5�;�i`�+k��_{�L�eRS� K���R��~��Q�d4��~)Nn�"���JYqrC�-��hb\.��$�>�U�ap`�{�2��k�?�ծ� �)enrI���Е��<���r4?"i��*0]n�����Ɛ�,#E`���E@�10��Q�Ф��@giM�2%�]Ȋpf����h���^JŔ��˳�`*�GLyIe�*��ƫ�H藺�ɡ8�u�R]$:�x���?{�[(��� _���ڷ�}s�0=U��ǭ��s).�d�<G�Eݽ}_��M���G��f1L�.�Q,�X^��]�����3��>�6��t*���j�<�X�ǝ[��7܄'?��x�&mY�pt�K���� ��,�^��~��f�� " M�� 

*D�QIbb���EM41F�H�X#�EE{A#��A����z۹��}�������$�3�0s�=g�����������}�� �"�9u���K���ީ/4�g��Vo�ß����a:*������4&�M���I�Y�V{U�ϣ��q�����3X�r�?�y�W\y�l���/��[����:1����|��w�r�8%�%� 5A�xa=�:�I�)-�w&r��g���$�2io"�xc,��J!=��.fX�&coBf�	�Muۍ�񌁒(�,���F���Y4�גk	3�
[�Tj���ԝ[�?13l ��筈iES�Gs��]���4�����%�qx�J)�� 5������Ç�~.�X��<kX�n�����~r���`�T����)Y��z>��L{buM�uh������$�%��s��L��bN��H�ш2��� �逅=�<�)z�Z�O%
=��4�n�`��r���b��+�f�$��o5V,��������!�.J�q��ڭb�D��O����Bs�읙Î=Sز}6oݍ�1[o���˱Y"����Q�Q)�3ѧB�2I�sU�+�!r�[�F�����sQ�!�A�}����I,V/�h�p�=#�TNY���/�(�I"�V�:z��ا���_���Ld3���?���_�� n�{:A}��B~���J�)+b��E�/�
m�`<�S�E�.�PR�/�TB,y٧�Ub�Ӽ��Q��������������n�v�I�Y�W�36%B�k.B�xC`c�;ҟɖQR7��R�9�8�w���Ȣ����9|������À�i�R�<��t��Uݰ+ƙR0鶲t4U�Ѥ��f��r��x�_����:q�>���B��/�|�j�����7s�%�[E�D��zﱷYD��0�}�M%G>�mK��5XGZ���ѬF`�� �_�|L��W͏�襴���10͡H6����i��rO22.�*�)���M,����c�sL��M�ټ-��j)�LQ�&s���}!H>jg3]�#ƔmTń�s���O�Eg�(�b|��퇠3	�n���߮�}�팀�[.:U~��n>������c:�l#��"H�6`� �`��]�畱H��6�j�"��=D⮥��]��yZ3��gpk������i�g�w�<�
�VJ@P1K&j��B1,���P��c�W�s&�W�3+�ys�q�j�Q�D�Z��&+2F�zP�q�ǚ�M�Y��-��j��F�H��
�A���.�rg���!��"��,k�	c|�9|�^��Eu�D���	���m���$����1��vAgr澛ϡH��R�2�� S&b�+�U(���DE����DB�UD<��Cb��@��;%�4�sLci�3�v�Xܵ>	g]�a3eS��4
�.��W���8:TLn-����(�{=4ՕWG�,��ZD�wg"�U=�Ce3S�޹Z��J��n���L�&�z��,��Eɩt�Jy���R���Ǎ15Yg2��PL������͇�S��

c#�~��\L�ؓb�F�=�<�X����I��G`�)/�)��Y0(	 �bY��/��i�)%x}q��(äE��.������
ڭ����w�Z��-gc�	e2���9|�K?�M�?��B�U�_3�3^x.�����W��߰���b�6��	�F�����3{�w�&;p�+��+ޏ��?L-)�!���ᾍਣ����M�db�\���[elN��"�Z��Z�o�B�|zv;�N!~���sL��k����p����/:u�Pz�-!%=��|7L_�|���RL������[w L�`|�
jU1�`�%cj`O��".���C�$�AU:+=���J�sʉ"������KAԿ;>��l�|�2}1��N���r2[Օ*v x��5�OF��b37�q m!�*ꟳ1NƦ�6��H��l�S�����L3�YL����b�������3+��k1�
��m����}ۥ� �Ƈ�ػ�Łˀ�� )t����_�߿m�!UG�4*g1�4G�V3���g��3&��֯%N���)�OT,^ӵ'&M�E9\�FY��C��*^�*�8������~��a��Pf�fRri�)d�0�f����P��"�>G�xA*@H��+r��~�A��a�ƒ�����P2D,��ї�-GhP�$6M2�G�Y=�$�6�?o	Q��Zx��zz6���ܠx��3M,��Т��$������x�mY�h����+Jx�/��g��M����l��i|��_a���,`������Fi'6��=Yt�
�O�1[~���bH��A�r$��-0M��3_�s2�������_W�!5��
�:��}��2���h&�_\:�]z�����h��u����p��d���_q�9� T��K#�^�� �U�ۈ��UXh��f#�x�ӫ__��j�p��RPg	�a�3D�ܤ,v/�!��?\"
�l�k>-8�-��o� fB�o�v��*Q�%�k�(`Ft�k����'�Õ����y�8��aA�����O��š,cf8�h��i�9��!lu�������&����g�i�����=Sh��������&��U&���}Ŵ�1%0�ں#fL+U��J�Bal#c�x~��_Cm��)��'yӠC`:��2�L�?=����5�+/��7o܃�]qx|��,�;���ůD-��m�l>��W�{�bn�/��#cc
�:�(�Y���䂪iT"��z�	x0�#yH�`�������vЮ�aОA)�ǉG��?��"���N	�}[����/������a���X��a����SzM:����Z���QF��SY�rUd�ː�N [�bH6���F,h�å&%��5�L��.Ha�oꒉ�.�`�:��(�Ʌ7�[�%��A`�A�mS�pb�֪�z^���IVq����O�o��t�φ�S�-U�n ��#aD�+c0r�a/�=VQ���ΏQ��w&���|hƬ����
�����bw����U���x�4P+����Gw�[�J^��`ҽ�xVz�z	�
����:[���#�T����5�}� �x
�`W����
D��k������P-;0�W`*3�XH2�؇m�{z��1��cJY&+^�*2�#�ӹ[f(��Q�/��L�^rv�9�-5I���86�a!�.�!RD��cq��XӁ��q�)+��1��@nb��*��AW]M	e6��@���'D?	L�Wd�aITM����!�<��C����I�`���\��5R�㯹{�X�    IDAT.�߈���O1;�3+�j� �9b>�K�rBӹ����!���kp�];�),Cu�����17���[ѝߊ�_�+?�A,go��n�����` I*%n�RY��/T���
���'�����XfN���GJ�R�>�fg$��g��˪�f�����g8h�t��Rl��
D
L�|�{�cמ93?:+G� ��|7޶�`c+V����N2��z���}��o����Z��
3�?��!0er����C��gFE,;�P�2?e<��B��1WJ�r儶���Z�{�45Hq���G�،�"����׈��	p١C+�ítU��Ic��z��X�E�@{�Lű8�����숥��k�9K�����Ϙ���F�R6�Q�4���.�A���<����8bu:�=����>�=�K�y#���۰��E~d_�%�aZ��EQ n��^�4ߣ�'��Y�3g���� !����ƭ�#RD�%o�`Bm�T�
�x��0K�������_1��u��uH!_��3t���Ig"�C�O�b��%�]>y_Ȍ�UV�2�����G�w�V*;�u}H̏%�V'U(+��c�]�����r�Y��9�V�I�ek'�0�/x�"A]����v��=(�[8`e�;�d���gI��ޙ�w@3 6O��Ǹ��)�R�����0׋��G�{J��y�B�)	��`�����覥3N=X��������!E�4*�=ݫx�x�w�[<6F�O�o˳"�)����dJ���$ ]�}[��Q�-5��6�[_s
�:e=*�kn%��?��x�>��Y���)o�:ڷ+I���x�E��Y�\w\Д�P�4p�����",��WЗY�,tݻ	x�_~��E���Q�)Q���:q(-T���.*�F��v�\1�go+Q!Y�'�-���Ӏ���c�S��1�#��Hy��h���h�|�=��H�K�R=�bSj��!JE��f0�+� �9U����B�7)hF~1�1"�����-����E�K�4`�Ӵ2��>c�X�-)7���8�� ��tc�:��q�+O�良L�n|��_���v0=u�9�(0�{+��Wp��07ߕJwmlT�V>�OŀB]j�{aOA��F*�2O�u���A"� ��r�9Mҽy��8��5��w���*�!�-p�V��
�{xa��L:����~�T����G(g��VmzO�JL��AQ����T�A[�Zx|�,��"�)m���Ջ�or�d�)��B>�&K�h����1Q4��U�!@�FwOp�H��ֻU��8�ʿF��X:�"<�@M�;)���q0Ѹ�,�T��*�X>'p��6'�ό.�y�'^�s'��&��&�/#{E6&I���0�|*�h'�"����DO��'Β$���&$�Cm��Z"�����xb�����ϪΞ�@29�"Bbd�S%nb7�(�p͈+$��kJ�s ㊔�7���2��c���d��	X0H��� Ӱ���T��͊�*L�bɞ�tOsy��3H�1]� 5RA��ݶ>��\��)����4�;���BDidje���<:z{��şߛ�)���c:=��BC�j&Ǒ���Xޛ��
^<Z�1�`Hg?���C�D��G*cc>����/�m��~��L�B��9��H���j�����{$i~�G��~z(!l7Q)gP���zE���w��FD�A�i������ �(��"y/�h/�aj�f��m8����s�}F�z��H�	��T���%�(�9�\R�;6oF)�C1Ͼ1�� K��&*�GDJ�N�1�����q�w���j������r*o�1�7�=v�c��e�ӳ���1�.�}���;~w�N�#˗��t:�()�4e���B���X&5L�5S��u�vɮh�"VA����>��-M�R>����YqI�_A��,��.%z����3�����Š�
����Ϧ��zDEa��9Д).�ir���Y��4�9X4���$�@��<g4���gI���1� #��v}a\L�k,��8�ު��2x���G@�Wrs l�����q�nƖ�}���BU�k�Q�QS����]�8F=�10�X5u��V�Y�� ��L���
����s2�F����5�hy�#��)O���&����*c�%af��K5�B�Z�����H�H��M��?qk���9�{JE��KX�oY����/Q�|I��$V^�y.rx+D{��1���ءx/~%�Gu�5l�N��<kÄ�wi7N�K<v���{� ��cm|�S���]!:uù���R�M(*L��̓*��\C�D,�SŒw�"�>& �+��@-7��@���~1v�u���ܗ�wU"--�s~�EW���+L�+�N���%��������Ȑ��!ݧ��D�ؗNA@�y���=/{�~�-^�)<���o~�z<�i�>{���CQ]�RЗ�^���ږf&BC���.��J��'��9g���L�ASr�<�C�ͳyd�+Q�HdYt�#_Z���?����p���j+�=$�aaɈ��c��#L�F�X=�b�%�i_\y92���dL��Xa=���Ō�����x���2.f�����# 7`JW_55���,�2Ts9�1ݻy�a/L�ǔ��@�^������G�2��,�(�)���F�����?�F��1�7޳K�M{P-ep����b4�	��[��䕸�M"����ز	tdF�V�z�U}��<���S2h��j�����+���8J-ȸ���<�aޘHv(��̡0�ƉG�ƥo��V�#E�{��5�k���9��+5��*���֍�Ǯ�A�G1Qɡ��@��B�1��h�.u��e�e?���ظi�.�,��2��nnc^E�C��h�#�cj�*!ъ�2��OaK�U2*$ɐ��3��{U����Klbv��;��imTu� l�xܭ��
H��/��2;Le��F3��e��>���fuNi:�r��̶�k�B�j? $�F2au���R� �1�<S8�P��S�����7�3�m����֭ͅ9�&����z�un�K�R9��ukp�,��jZ�V &���(������NM���CS�D�;�Ъ5�}h ��Uk�V�Rh��L��B@0��N�0�7�Ve�wK?�y��b�V�J�䨱�c
xh@��PdoS��ΞY��b��J~�ZBq|�BF�����+}fLd�Ĉ�)�,͏RLʔK�O�!3RE�� 1�B���O-��4���v)���ڐo��)c�4�d��;t�^��!����yY�G^"D�9��}�ᆛR%��&j:v�b<�O������Җ4�m�Ŀ�����Ȗ�A�cor�i/`j���㨃Fq������A��������U��j���e 4B�ھ#Ŋ��=2Nq��8r3i�������d �=�?܃؈��v*V�3M�t�d������1���A���k�<>bLY!�+�[��3���L��&Q��`H���|�%��V�d�Ζ����@�����Eߜc���S���`	;�	��Z�X�	�W����'�"y�B��MD��i�O+	�0��'��d ed\�F$���s�|��{\�H��IW�L+v���~HR8�Fs蚷��� o$�ث�j���'Z�}�d�n�M�RB�����֕���x���D%�4�8j�N5����q|���m]��@����t�7o
����2 蟖Y�5Z��]��P��a��,��\7lV|vl!E���z7w�b��6E���Ibk����*g��� �3�=���f.�Y?S����������UvUש&��p�Jt��sSi4O�G���;{�E���/E����׏[c|��D-;_"O�d�9^d�Q�8���^}:^𜵨e�GM��d��Cຟ?��~�טiЦ<�P�65jL:_k�����r|��F�:�q~8^���>\�V.RL�-�����E��b�������w1��U�E*�%E1/�' �c�{����6��؟����RU@��ϰiG��}����^gV��_���8����<3k%t���� �.�}��F��Q ��R�U�1���.Ϧ*!��c�d�#)f�x,pړ{�W]|)6��Q[�BM����!C�H�b���'�v�z�c�$��J�5�cA�� �8�4	L�+�F��J�i>/��=��=�9�R�R4 �?�V��_�%+ �U7�A���N��497��D������������b�t�=���BI�T���&�ˀH��z>��\�);�Xy`᱇!]y��L����<�w���C���g'�����'��w��xǛ�G�ӻ6�]����,�4>�Gw�-zv��OP�I*��3 �z-.���<���('�X��ﴀ�Ⱦ��Z��Hy�8�ux�_�
�V(0%c���j��h�N�|�&F�l4��^���؀��@�cM�+�ʊ��+q�
�`w��;q���b�L�\I�SgOCt��oV�,H'��b	�:%jOR�40��v� ��u;v��';�"�x-�'I��ʓ��,��	ǆ9��ŲW��6�x0�b�k�DL�\J�i���P�!Y�Άt��� f.��]��r캣Y�z`E���fZ�`��V���i���1J��>jb��A���~Fa9|Hp4�+N*M;h���%����NL	��x�5-%+č+{����?�N_F�m����1�
J%��rЫ�Q�������L�Ƙ�gfі�-=mB�B�d.��b��]M���4���DƴV��Vn�o�P�AU�a)� ��q1m�tq�Q�:^C�@�$5lRP����3�-����D�r��H���2X�A�Ta��K ����ư�A�}���2��D� .��u1�w�1���+r��߾G�/I/������_�?�	�.U]��Y�W��}��o|�_;.�Y�3�ǯ�>��㻑��Du�*}�"[k70�c���q��*���G�j�r��J��"���!fg�h��h4ۘ�[�޽�صk7�g0dpe!�j�*8gCj��H�V.�~��Ӟ�~��9�ܽ;wm��-Obͪ�x�K_����!�5�({j�7���k�ٹy}�\p���g�ܷ1���_��gp����0x��Ӿ<��0�����߬�I�N�M=cz�ޣ	���C	)f�bUB�Ȥ��$��KVRqN䈞F2@���G��1��x�-���T+�1�E�y�ʗ:�G�ؿIA،�"C6�7�9�)0[l��b��Z�s��kH����uo���3U�¿��A-��y���[_s6�F��ܙGv ����q�����E��a��uu^�I&u�=:����R7zs�H�M����d��C��~LcV՜��r�F猺�s���v+�D�����#:�
�Qm�TX�{I�nc�\)$癵E�������$O�{ί�h�g�_��f�$��E0s(�S#��<�����s���,%���"Xo�H�-R�c����i����ngak�t'�?�ꢳq�!�������zZl�x���\�C���]�f��ry-�Gս�k����X�Xq�n�e(�7�0l��6ܤ:��
��5&$_1���/.�#K���W��i��Т�>�x��?A��i'�D/}�*��"O	���R ��|WMmɬR��`�z<�;^w*�8a� S�^#T2'nK��4����ş|i�/�/��N+c��་ߏ�3y�FנX����=�Y+�`���c����.�Kd�h��ōjSZ�5��i*�M�8$E'�gʨ�r&�p����,z�HE[��L��2*�g>!D�Y�x+�(e3�Zb�Ԭ�ud[�8گ��bd�,fu�����bƔ���.r�$0%�f^ K�`�ǘ�i1��,�ו\kH�Ό2��:��<��'sL	Lo�g� �7�`z�iG�o�@�)�]���O��M��ibb�jc#Ru�<�	g�2�a�f�ny����1"�N7V6Ƀ� �8��y�7�}�i�����1q�b�"�A}n��^�38��u���_�Փ�do��|�SWc�óh�
�O�a���1���٧����DcJ?��ۃ��'k@�!C��!>����C[H�k<��yP�䆉�f�̙�6:0|̋1��[(v�ɭg�cV��B7��()��.��ɗ����Yg=XԭP�mI�T$@J�XL�%�ɬ,L��&;�`�VB���3Lv)o6�T63�e�ߗ���IYuMgHZ��!����W�$����c�W��+V��[��wG%�:�U�^\�V���:6���y��e�Y�e�dG-,�S��'���٭�Q�LY_:bH��E�05k�(������80�
��%[��J�����Ja'�<�Fd�9����`���=@)�NKPm��Y%0��1��}>?I��4
Ôӽ��ͷ���;7ZCab�-$1i��	V�ٓF��h�;SGg�!c�ҥ� SJyu`�>���i=c�)����\S܁S�)���L2˔��p�C�u��.��&�]\r�I��e�Kŏ1��y��޻�Nؓ}R,�˧Qȥ09^�<�=!���n��/�~��'���@�ʹ{4_�m-`z�t�����K��`�R^&��ܱs/����d`�>���ض}'vOM��h���ju�l��nvd?)��q/+[*��r�դ��+�jc##�ȇ�:h���g6Ť����z9�y��X69&��O��~w�.|�G�K�?�u���c��0�Z�읟�M��q1�+V
cJ���c=�:k*M���%qRWuM
Dz� ���9��K�����]mq��=��C�d��m�z�"_�X/-9�t�]�Se<����+-f*bw�4�Ѽ��JHʹ��	�To��l����^���@���W���0�J;��+��x(�/��1�������#ߝ���K.x	^������4�Ô��]�sb�����b�W�07����LK1�}�|�4+$xҢ�JS���|�~�0vۤӢ��u��F-�)�s�fzz����5g`�%�Z`0W}o_t5վr-&�?G)��R�x���xT� B���:fD��z�A?_̼� G�-fn��b��n9�=�r����$���h�)��Rd�ڳ(�x�����~!�8hcJ���b>!s�Ƿ���o����Q�m�FE:Io-<Z�O����A~��҈����{v��w��u�V�I���+��-�)�U��D��U������ş%�����z9�8@�skQ�=��Y*���JsNm3�S*�*�^L�t;3�wl�w���	`�3�5����R�d���&	d}9F_����)�.=�O�ν�}�6W�^�\U�@�L^�<�?.�W�ϓR�A�.�φ�aC0Eݩ�
��A&�BuC�ir��5?�FLɘ��?SG��)�ft##
L�HQ�g�P��� (fU��o�� �t^�C��0S,�k��b`J���aL�\V"K�����T[�K� �"����60lMK��_��|����K��Y���
Ș����m���\���L�TL�ӎ���t>Ʋ)�'���.>q�7��̵019��e�{]���.����r!�/{���gF�<�M�v���c��i<��V<��<�y�X��ؓ��"�2*c�
��L幹i4f������^�K��j��,E�������*�}p}��Nab���r���k8�Ykp��X�jUpm�	�iar����2k��x�f�˾�[���'�*�櫀l��Y������¤[�m���ťT�{̵���u���	.z���j�S��T����y�O���*e�ـ�H��P�lҘ"�犌O}�g���}2_ИM��GS C&F���6;1�4�����;Au��7#�ښ�/V�@z��F�Y�IFm+�L�.]�p�%@vM��ћӳ�_�)2f%���%�k�$����ҟ�7��2����z�n�dQV%3� ;K������7F�.��=��9��Ѹ��|���h���:H�Q�q�iY���dL@�'���;�IW�1���Y�nQ�Q� �r��}5Ǖ7%h�JyS���9�O@#^    IDAT��3h�ѷ0Qà�A(&j>���+�S���ҹy��3�"(搟T`�Ϫ;�2��YuS̏��7���$`��4C� �i����i]�Z58��o#��������X���p���\�� ��A+�p�� n���'��;xlS��o����7�0�s3͝8d������5��L�Zܓ[���U_�v�E���D3�dJC��u�s1������it�lQȁ�D�X.�ɬ�.3&�����Jd��(�銹�t���z�֮]��?L~ONN�<���w>�w�s?����#��_�|�5�_L�ՁK��2aLC�bb�**5�����Ė>0����k$m���/��Q��;����곎Y�d��\="�G�%�ۋ��',����I�W��P��$#�@%���l�`��ь� �&����K��v���[zea&����~)�TڌfY�֮�I���RF.�bv������E5���j|Ց+�`����38�������XS�-��X9���Rhr����o��"�ҥ	�Z�s�����e�/j,)|H�I'd}=iU07r�L��row���/��S��0��Tzq��/���v��{*�sG��ͻ�z��/_�������~������gb��颳+���O4�y��  |��Y(�������K
v��Z��n��>�I>��{��r��찟?��w"�W�y�=���'@�r6��g`�� 6@ɿ��;��~����,*�T�e��ДX�5����c�g��+��9X�>QyP�#���R�]r����nn�����|/������w��#ZˉWڗr��g��r�`l=�L#�l�J�DB�+�S�~�δ����ׂ��J�D�풱�vM�X����q@�w�?T,��whC�F*���>N`���a�B��*d藐e��)�"�s��Eɢ�)�U�}����Cno���W��4_�t�e���K75UW��2.��͢EuجSu�u�T\qM*��z�P�DG^Jy�NϠ9���:.f�����c���XH�)h�������	�/VP�T��_��ڸ!i����̝h:;lNc4]�%�<o>��s)��l��>�U<�m�|g������c4����<ⓟ�n��Q4�=�NT16^�!���К�h1�1�����D}�A���)VRi�1Y�a4�0�C�m��?�%�v�C�Rj��#[.#]�bl���#Hes�!��yt�wc$��>g.}ۅX��$2�{L��+�}Π���F^_6�� ��xe����b��c8��58�GbbD���{����?�%��z�)8��g�2��Ǯ�oފkr���$Nܨ$)O�{+����w��\0a/�I6d_�S����J��0
8���=���j�4�ZLt[:0K{�MQ�b��2����n��O�	�WIcFQ���(��؝R�\�NȜ5ő<J���2��J9�Ħ�̽7KÎ'}L�	L|��N�����~�sk�X��@�EDze@�3J�[4���""�Ϭ�}^��_w�T�r���=��b�8��M��G��'r�>]���h���rQ��
	���qםy}N�����:l�.�G6�r�,R^���1��h`��"#L�29q�W�w�A�ϚJ�s+��M�ZE�!�i4CU����1-�`�(h*c�9�4I�2";��tX�+�2�*7���g�#�%[��Dwv!��N(�inr��8d�V
n�����wʘ�.`�l�#��/s�	��ϐ{���@�1[��}aR#N�!�]@�7�s�8v��؇.�tZ-�}�&�;Ib�L�����=���n@�- �)�Z-ۈ�4���ٻ��.�o�q�G�vyZ�h������|��3U�l�)�yٌ߲:������6vO��ɭӸ��m����K(W*ƈ��NZ0�]��&�� ��J�6��a���c�br��Sعkv��#��kV���}VI��<砶�zX1QñG�c]�� k�Rm���]���B�_�ĪU��h�N�R���XXms�6Wb��&�%�[�L���j�'���h+/>���SO<���JGW[$��ī��/JD]�F��q�Cb��ĪK�|���$���আ;
8]�!�����I�,QʳD�㥽w�5���'��C��׀�����G��t��
A��)9�1)=�kL#h���G�w^�*<�����E?#fL�.���Ӯ:p�nǗ��+�O#LU�*H�Н�"������L0e�ZQ@�{OE�l#��ŒO��E��I���2�zG��\O�?v �緂ac�#�d/�jz-qJڍ���g��@z������1B<��)�+���E�v3e�j�K�]������*�đ��%# �粌�&Xw��7�L�.�_=#6�k�1�Qδq�!���sO�I���%#��U�Љ��M\��_��7ݏ�����'����=�1_]��7~_đ8੠1*d%&ĳߓ���Xf�@%��1���*�=	���3���B�[B�=��ދ���[�����%
2�o��s�')�D����J>�rY���%'0�ug�z���i8��"7V% l�,����r�(~d}��	��>�e����s��Gw��}�ݬ W[�t�$�)G'ə)�1��\~/YT�P�{Dw��_[S�.��Ibx8�\�*�������b�)������Q�����Pr�P��� C�V�kcƴ/��li!�Ơ�`ڨσ����Q���x�ɣS�d��ธZ��A��=On� �"W(%�)g����L�� &JL�1uc7Sq�H�Z4�b"��7��x\��0���[���]�G�ϡ�O�S���]|F� �<��]�[o}�v�RccEd�]���x�3��O�}N8� T�fE�ĺ�b��Bs�[�܆����ȓh�@)H��O��E�KP����y�vT3�v�Ax�_]���e�4����?��M0�iR��C63@�5���m����q��U��GߏC6�+�43�������Ƶߓ��>�(���=�_���-����}���)�-!�6C�N�L�	L)�]�:�ʮy@�%(m�er�[��:u/���� M��gȸ��� f��XO	FR���OV.�ꫝ�d�2dh�ڬFV�2����:r�d��ɔ���LQO͓ܞI�W&!v�9uZ��L�h�E�n�$0�\+���1���gN���45��mdO����y�Ku�yo��&���zht�_�ɳ���\4��X�L]��Е�,(�3{�DG�|��u�.���g�d�JqQ"_�V�1�17'@�U�Ō��8 v)W|R�C�8�ղ S���ԛ�i��(Y�R�Z왠��l�Iy�.������� pO��i~4�����S�1͎V�O-�QP/��L)�%cڛ��md� ��א�����M%R���qU]I��ݖ�E.��x�G἗��5+�Y�� `)QTwP��q���،�|�'ش}�l#�1�GRXqn,�bvj���8pe_��c�d
9��� ��z�	L��D�[�%�v t�@3�޸_��:�t��@��l��b�"�����K�_}΄��^��oy��8��e2�\֠��HBuhu��Ǳp9�KVa%���L��Y��y���m��X��jdĜ�n��~��4�RL�����R��{!H����TP㙆'��ߵ���09'Y�7_w�]�t,�^s`��&nq�ޓ>e�����N0�����-arĝWю��h�@d��-�����X�,�^���@�Rgg>���̝<q��l�?ǅg�&fJ��1ɼy$�8�IX�ϣ�ZeM�T�ð�Bsf'��i�����sĸp,�*%����#B(��7�>�/]��q�v̶RHF�O�-UDʙ��:��8"Y�S�4[Z�d���		�V{1U]gM���2PI�]%�ӂ�����DR����"D�m^ڦ�o�R�{�����%���T�]K��0+2}�ˋ<�4Q�(j�T�����30Ձ9�
�,��N��;��	�LTsХ�)J;�C�X9^���=��y8puJ���#�.��2��Q���?�k��+���,ZCI��EyG���MF���=�o�&'*:�8G̠}6���G#�Cl0-���̳��.�|�`��b���G�,�����Xm9R��������`�փI����@�8�b?#\ǲ�8.�K?�&�y�[���\t*^|��H�ɵ")�0�
���1EN��j���G=�<�S��yV��{/2ߋ8��-C�wѻ1�Cat5�ժ��c�X*g�X�����[�<�&�^{tJ�h\䷳ &E�lFSe�ȍ��EYgÁ�nvW^Ӧ�S�� �͌� (�*0%��"	��0D!�p:h������)��dk�h��SU�̤BSC"`��bڡ���5��@e��H�-ʔ ���SG�g�ٺ����C�ic/��x�Y�ş]p���D�o�Sz���V|����mu�:�����7�+��7������s��ͷ>�f��Bn�ɉƪ������^W�$��nT1 *�A6�n�����E�1�����m�-ܲq+��{�w���z���^�,��3����)�,c�6�߷x��/�� �Ԑ/�Q��IQ�ۉ��-(�zX>��Y/y.y�9X>�R��f�������E���S��K��Nl8p�8iN��˿~��ѭ#���8���U1�p�z����R�ֶѥ��ٽHj���$�GŲ;Kt����hH�W�2��>�jQJLi&kX6���-+X쯓���F�@A�搩��P6WV�w�Y�qa�`��T^:��x� ���N��[$��H*���,u��!/t30�I�G	�m|I #�Ke�=Ӫꄧ��2K�`�
+�#���=Z�K�Q	���*Җ��-2��"m	���o��%�{��k���<{*��Aʘ�lq�%C�>��=�	�v���u�{i՜;���dS�ajI.���1���%) p&h�l��i���"�i�����?e��!:A�)��I'g��L3��v`�
��G��E��S�?F�4-��x?�����ҵ�s\�,{L��;W� ?��ZYS���nȺ` �g��Jy��9��2'�&:�W�:i�"ɲ$���{O���R>/��A��Ɗ<���8d�JL�s����k�s�7���b�lO��M�?��;[Heʨ��ӟ�P�i�Y���.��Vf��>������Wŀ��Si����8\Rm ���:p������g���[D���͉��ES)��<�p�p�YǠBK K(�2}���m�l��t�� ����|7߾�^I�)Y-SJ";�c���{�#��?Z?���.��5�ɹ�V��=��*q�k�O�"	�M$�Qd�f.�D;�9���(&�d��ů(�G�>fM"X��,����֨_>�;�}�Z��~Q��wB��@�Q��u���y��N�Ҽ_Q�GtWո�=�_A������iT��^S�&��;M,L�B�Wǡ��x�sO�Y34�\s�'Pi��M;����\sݯ�iw��$�BM�z�f���,���0$	�#Z��'�*�q��IQ��Q�2���W����˧/������=��gڼ�����G��ڜ���m�2"�M���h5:�L�KI�R��nD�Ì}"`1in&�X�SJ�T�^�_�~�Zi���n#�'�g�z,N9aj��1���TC�k�,���ދo|�l��_� [E�PQ���%�I?�g�{BbW)��r�n[�Q����bLa� a��?����[Rhs�K_��4�K3v#$$�qv����ϱ�0��c��'Mѡ��b�֢�B�'�zLUE��2lc8lb��}ѩxɱ�Mʫ����#O���;7b��EHu�.�7����k^ź6��:���e҇�-���0R-�Y�<�L��ا⺹�.x�{�ПDq|-
�)t�,\�ic��ss�ޏ��G�b=ɖS��z�K����ˢ����<Z3�h7Z谧�X�SSJyY��)��E\���L�6���&�2d\�d�e-�Y���
�5�i3h����]�KecLsږH)��-��J"I��~L�zTN�(�P�)Z3�6���?~��ki���������_،O�L�� /?�0����c$G{� 7��S��n�e� �J~�}��q���������F�cD�c�g\.J�4��Zg22�e@����~�gx�ɽع{��:2�j�6^t����;^�u�9O���ܿxץ���Gg1J�c*Ւ�I�u�!�=�@�vҳq��`ղ�,Z�`2�7��N���B�\�Yg��C����6�?����~����d
 �"��2&�'}Q<�(�BR�V�i�<�(�����I������J��<��X��TAZ܋�$N�-9N&�9�<2r��ep7�]eW��'���^�;�L'nq��dXS����=M���B�(@GG�5pӘ���,��03�u�>c�v�@IX���$Pw��wd����C's��@#�wȐ�(iU���@(V��W�aˉ���#jīfv��Ǖ%V��G6�s0��Yr%m�L~n#���>�O+�̝A�	p����C�r�xH؉�C�H�TY{�,�u���ns�d��s����b�(ϧ5�@�#������dɥ�͋%>�p@l�ŵP���֥����zLj~��g�f[��(��!;V� ���-=>�䚜Q�!�]L`�'����ϰ���^��}��"��N+D~h�e^�P�_�5�9�p`�qI\8���s��4�j�la�m�ߚC�9�L��젇����0HQ�L�M�rH�*��F���� �h����%��46fDʻaU�������Gv2��eLJ�]�O��RS��̞��&p��n�_���}�TN��-�#�t��?�g=g1�םw2.x�sP�0It���u�{����d�c�F��O�'�L����܎v��k����
���H<e�O�|�(�+��-�)���먇]{	��6!���L ���hIޙSu�L΢�Ϫ��ti�����������`MV;��וqO5Q���6?�n}���=�{��){��ԫa�K\ɸ1��H��=��f��Y�R�x�Б���Z���Ɇ�>��j�e/d{s�w,���;�~���U���<U���̴�[�Ʒ��;�p�Ch
9u8]��}��5�{j�N"]�qq�Ba5�28j�hlud�����f��d�������{c�ݞ��t���O�m�=3?k�z��F��EZYQ�7~v2�)�u�Lcg��j�|rͱ���k8U�`}���t�� 5�#`!pa��i��t�H��a֌�����ӟ4�L(sk�v�荡�RƐG�����ߌ\v͑A-c J�	NY�P#5]y4�b��&����"`*�����-����/'Z�fhwP�z�(0�n-��� g!��h.远9�׳萘s��X-:8 _Rղ���'�BT;���u0&~$���눕�oRo2wW�pT݈��R�&�W�x�O��ǭ�q1
J����/�W|�j�>h��4b�Fo��Jsp,C�=�����[X����V��O�8�����y���/���ZX�|mr�B�K��{�E���~�)�@����jf��Zcn�~FS��4`��<�aL�!��*��7���K`�f�U��t��T��~z(�O�`�}.��)��r퇡 S�y<��d\�d*
L���`�=A����){L9�1_��X�
�։#ZT���p� S�t��fA2�.R����e�=~�d$�TOW�5�C�an��V|�����3�e�8���7�J�Eqݼ��O��5���)�s�N?�h����c���\�8]\�M=�wy��w4��B�^IL����o�����}p;�g:�,�Mu1V���=��?��	`�x�.��͢;(H�42RF&��������⸣�b�
i4V��d�4�1`�'��cK�f�S&t�,>�ş�Ms�G���D?��t9�U�� �fC�z�6Z�ut�2�G�Qeɸ�����t=#��4��a�;�Tj�i��#�����5���(ݒ��H�\6'=r҄Oc�n��٤����� �c*���|��l�����P����    IDAT~s������)����b����\��,�g���T��|��X�2JEe�y�%�~JM9ϖ`�2^&/�$�4�W��
�ܜGl��	.��L5��2dO���x#��zs,N���"�k�'+FP.G�{�X�������I�"	�U���P)�ʏ��=�fr"�W|��UX2�*�R#�x[�aԤw�F2�IC��0���ł�n�_�ٖ�W���w�b)��M�܉�.���C���Ȣ3��T���d/������S�c:L����q�!0|ε*��
�0��\��D}o���2�>z�tgt\L�� _���bY��*��L\k��M�cJƴ��\]S��V�zPj���k}Ò����G�l2;��!g�� n7ќ�A�l�>����L��7yd��SOi6TD.��~l$L��UQ���m�1l���~\���:�����]��n]{�Kh�h��G7�����6�˓Hg
�*��##=���M7=���^t�3��o��]��q����U�>
m���KN�����1���p/Z�V�]�B�"�G��'0�R�<Mԥ(�E<���B�q%4����"�$�愙0K�[��>�[�;#�+Q�� iI�U�F�OZ5Ê�Q�bC�5��Qe�z����Ǭ��ɱ��"DQ�l\`J&�F�8J���9��G���K�W�8�m%ѓ�	���V�g��0�,��{.����c{���p8.:��8����M�,�g� ��7��$>����M4zyre3Y��Ed�i����9<��)�l	���� �Ә�y��G�������c�<׻�RZ_#
�4�J����C�
o?��IsD[֋���VEUe�T������S
��j�ǁ�zW�߅�OSz�~Ү��ɚ��XV^r�x�+O�aFPΘ�_
���$�[���\���N|������w��I��/ Ȕ%�b>��/�	:Cզ���SOQ-���n��/n%?���3Z<��b����|���7�k�DaH��x��?Cgt}o*p�D���ƍhEY�W����D�ֳ׌�L) �˱W�)��/"���cL��Pr�T0#��ci��u���V�����&��~~�]E�������|���G����u]�^��^�MFT�8���ɏ��E O.a q����w�C��N��
�q������K�u��}HV]cc+7�����ȟ���L��9�1�q1P5�:Q������UN>�o��WӴ��%�{a��|�1~t�O���B={LggtN=y�<2���15�$V3YTY�^h`��tzȗ�2ǔ���xS7ړ3�\�U�;���Tj�)�)zM�=+��O�8��Se䓛:�+3�?��@`��/\�G�Ϣ��L�<>~�ո��e��D�����wֳQ�Z�i�h1[5�6�B��m�Ĳ��"�� ��/���#<���-:t�Q�1R�����s\���2�n�}�a�#Sh�8&��H�lG������s(��-y�i��M�D��������_��;�b��F._E���g�����O�Q��ð�p��m��M� ߀'(�Ŕt��0��U�1,JxBm���L���X��\'�^������ ¾�,�L���*UM��:f����h�1?�a�t�]�Z'+��D��=�k� ��}�k�5����s^�;��X�*T*�66.���4�`�'�Ƙ
K)	�&���62d�(!���(I^��P9�ψ�&�u)'1���8ϕ��L�-<����<�!ln�>0YMF�dk��'��L�+����$�V5Ub"��"����}d}Z���_���1��s��a)��ߙ�|^IP	�E&�lJ�<�iZ��6�����9>|�D����d�H�ZYS�7�����aZ�Ŕ��2�gJ�0�� ��47ZE?�.q��^` �/1�"sJ�Y��N�"�o�������LF�G�Բ^,Y��E�6��a}�6e�&�#e�#�"R\�k��q� oc�x3��Y��f��=���M9�J2�R�"�g@��lF��ڪk�E�R�
)�:��uTsM\t��q�A�b�XQ���@���<�����V�a���\��'����߈_�p'f��d2y�g��w'#�G�q݋��9Q��s�p��ar"����L1��݌ZrQ�Ei��Tc�lޅ���^ ~v���W���9��Mal�
�U�m�5+��k)`r���U���܋R�2C8M�g�\+��Z��P���M���qx�E�����T���4���7����ɯ'-��{�z�u�`@tJ�g27����W�W+��e|�:��~]y����{�K
��K%��9�W��@�&ɑ�������kG����X�jr��E,��y~v@s��<��0��/|�?� ���¥�D��j1Yd�ϣ�׾�K���{�ywAa�W�-V��K���Z��SE�n&�0z#4�2��I��m�<*�y"�`�� g�/O����dV��M�ш������&�g# �e�V�P6���������K��7��N��K�6�s��@�U����(��g0�ԑC��^qƉx�K���Ie���\�.��� f�4p���Õ��%���ER%�<r����&��j.��B��)2'9��d�F�I�f��ϖ��6�n�)b����5�^[���y��1��r�QQCrSW��3��^�il�Y�HG$��O���e�p�ϯl��_�=�p߻L3̋ҒS�ˣ�61��ᬓ��O9+�5l��]����"��j`�*�2����e2�̅��N�P��QGE�Ԁ���62A�����y�r��4�f����ݍ�^�4z�J��B>�Ǌ�#z_�^��や�����Ѩ@��9��p\�)���B��C��1ͣB�I�1�;�c�/ Mp(sLI6h!R�j�\P5����+/�孶��9�U��EaL�,$�9klR`�q5L�a�R�ڈ�6���J&-�Ě��?y]MŶAq��[:sM��5������0�����m�e_�o�A1������i��ۧ��+����y���{�*\�Æ�e�x�N�W��4k���Z�7���!p����/]�G6��IR�>�j<����w�V�2�u�ʻ���|�
l|hZ]�EMcٲ��)�v���4{�r9�H�5[��W+�j�
+9.�h����Ǖ��~q��id0L��+Q��5g�M��uD���h-L���b�d�AGf�*� �YaM�˒$�uJ���{�Z��V�diO���poi�n���v
�����L�l�TLm��L�	8 N���@�1�N{Ff���M���l�)q�],�*�p�D(��].Vnr���TW�u�Eq�:K�p�߅�(��"
�2r�� .a^-!@#����|v~�^��8�R[���"Z�JJ�DЪV#u~%��<7��$ت)<`�蚑��9�E���FfW��H�N� Cj�頤B/ T��9%S'�-��Dcڰk�ଘ8��3��	aJ��9a���T,kʃ�մv�!��O&����S��St.��"8�"]�-?�Sd�٫��&�A�2:.&cJ�V��lN��sc��**k,Nu&	"�%�
#��NϢSo��d�˕V.G�R�S�
Spi��BJyS\��.s�	`�C��3Q��i�H2Ps����k�Z��%Z�h�g��9�t-�K��F�H�aJRI`�/Q�Sg�I@Ձ�L����hN��#�
9���K�ͣ��E�͋8���ϗ���1[���]{�ؓ۱g��� �\q�9��d�|�w�J
cE5�vo�r
k�L`��Q���~�\N⠿����8�3t$�L��h�h������x�H��Hgi��k*�T�4��d�*��M���٤DBU�P�N��U}�$����R���$Z$w�DO@�K�#�7�>�1�?xg_ָ��*=ߜ��߁�����$��~����5��-��͟Uc��,� u��y���N,M;�Y�bΔ>KYSY�>�2b���z��˩��M�<�5�)��Z9TQ���'�gp&:���,r�������>�x�X5�㔄�M���_).�ݳ�/�������7#�8�\�L^dr����:�D��hV�1 >�Zg�.�Y<���n�)jdz��m)��>��	
�8jg�K{��W7f��U(.��~��j���=5�n>�kE��ZDu�X�9�L�?��"�𜩋$��cY-�O<�>�<�(���s���1��,Sp,���B|�������{)�5�9�+�1I�O�g�0��s͗K7U�Kz#��P���������ӱ�ޫ�tG-bD,��
�!�4�����(+����L�|��þ&�4����$U4�N�N	@����ĀQ�.���p�@-fz
��6r�`,?��c�J���!�L7���)�zJtjfN�|�E)/Ġ]']1��$���x&l*w<K�頋R���X��k'1V-����|�oۦZ�+�!+��\Z���5䌙��@,q���%ڪ������e�1�h�)�"��S��0��S���<�j)2���4��Ѵh��z�̙�B8?3�F�,�S�U�S���X'f�4"Jɨ�2�CaL���Ӹ��y5?�?�XO�B�_ʘ��:FR��0����7?�˿|-�1�\f��O{�~�����o����=�Y�^w������Q����U�t3	�e�8�9<8�f����V�k0} �}�:<���n�`�:��^���b�$Gp+0�����Rއ� ��ąor���>j��{�zx�rö�`S�󘝭�R(b�>�8鸣�rY����X�����p͍�i��h��/�$������Ҵ&-Td��Y�;�SNx^y��X�|D���#@���l�tYd0����Tg�ǫ�z���Q�3��d�yW��魸��'���	N�z�Vƺ0Qv��	��(f{ȥ�8��8�ȃ�l�*,Z>�A�X@���� W�9�V�����=��d$A�#��3�ԖOM���wz�;����o��SsLf	��b��
��Ԝêd�Ұ#��17���^��:ݎ�KҕP�Ԅ3��z�{��J/�E�k���:3&�q���L�E�+�����r�"����b�YsWM��6�v��0�R���j��S��SC�@�X)}�w�`�;F��zT��@��Hz9KE��e�]��T̷�44���ʖ2qw�#c�������HSRhs��edmd�<W�2�dM5`
2�=,����1��v�նc��OI�IB(B/���HQQ�`��bA��^�}v� �(��# �� 	5!$!=��v{ߘs�k����/�s��k�����c�1Ǥ+/�h�N�ނ ���=t/s�%1C�x�f�*���<�S�g�$K�* &��� �g_zLh��au�Iy�	Y2�`�@��'i�V��Y�N��&V���i��4WhM �8��U��̒K-u�<G�$��w�RI�K��z���W�W��F1$��Gd��q��=I橈P���Q5��.�)��:&��G�����z����Ew�q�k��7�z^�V�ʄp^�R�sqIx��+��Zm4�4���<IV���E�����i�cq��9�@	ߛ�C���o�jB�������F&�&��I<&8Nue=䮗��*�51w�sM�t
W��C�c�|`�8;�������;�V�/ÕϤٷ5��I�$N6WV����?�{����kB"ֿHy�*k���N�[�(��@�[�Z�քVq������1���ĵH`̙���&+�U��@����-�pw|��c0gf֯����~^�/i"�3���;���}���$Vm�@'�G"߫s�S��e�LS	Ź�$4T���HK��~u���A"�zF�`s�Ys����+@I 2�L1ٜU�$gR˗�;L�A���'�v������T&>Ybd�[���9)�VRu��N� �*��[*�h5J�*�$��s޶8�Cq�{`�i�vN/,k���p{R���+�p�����U����IЉe���3�#>(�2�:bvFj�1`@n�mU��T�W�!d��->�rC�{6n�
��d�0�Fv������
ֲ叡	��
am�]o\�V��#��	_������Ҭ֦*h_��Wy[�����ql���a3�eJ���p�﫺���c�6Z�1!�:����&P�D,��ILן�%�m���K��I>)f��V�\�	V�Muzn��2�mK�kvQ�$ϐ�`fN�P�����w+|�䤓���>���|Ϊ�nJyi�E`�C4���#bL�b��)j�VHVLs�(�K>6!�R�)�}�f~��Jn"�Ʋ�����cE��
�V��n�L٣ڊs����zTE:G>�@�Z)o�c�i�"ΣҾG)���#�d2��BT`*-J�LY1%0���Z1-𶄢���"s���7q�b��2��N8b>���'ћ��@�{Y�����|w��.~��3p��{���&��`A��>�A�J��a�?���ڿ�d���s��ފ�W�a|�)��b:�b�á���>���t�.�ު��^�wWO / �J ���UG"RC�3��S��e�6�c�+�g_��U�їM�_�4��k��]�c ���%���ǰbm�HF�?�l�|V~F?��`��S�@���~��p�N�\y�a9�{ew��A0��� �Mn�y��VXLUx��	\s�
\yӃ/3��"��3�� �@`(e�"%d�]@\E��]w��SNZ���@���N=�,�s�r*��́Z��9ms��J�W'W�Dx��	\}��x����ED�/b�T���	4Y�q¤{ҿ@G����2{3
�eH�]`/M��!R�\�%��� �$/���Q2:�����d�(Y�F�������PB��̔�2�❋2BM�"�EubT*�MJ�H
HUM]��,��|yyz0�9t{�����k���bРĘ�>��$�h�b
�&#�NK�Ńӫץ�Ɋ)�	��9�:؜��K��I��z���L��xON81zr2�V�������-�6��^����}O�b�TL@"�R��(1?bŴ��RE*��|NzLY1�|P�
Sv<�3��{��{Ke�i����QÄ�h��[�U�c��"���]�xQC���2���E�N��^���*W�,q�3�,�ɢ�V����ie®��*g���&��|��5(H���:"��Y�ɹ(~�b3�����W�5bE������ë�^�I���4�4Y�r����gJ��j�"����Ӊ��L4b�NŬę��xL����䫄���S`��9�2�ׁ�D�U�TQ���Dr�=;�BrWMҬ�]�UFÆ!<���8�W���f�9�����tHswɭU��$p���S� K1 (������/��Z��Sˍ;�3�M������D̞��v���"<sM%L-��I���"I�i��ώ�� {���&j��&�C�����WNž�o��^٫���s��p�]��^^6���xO��Vo��͋z'���d��#@�ʔ�H�^���� �y��f]#��p�.|u�˃$����*4JŘ犄kI24�(X"-�L�4Z��g�R{��o������p,D��L��T���iRW�al�}Gh�"�~�GЬ�#�m���n;O�	��E��̩t�t�� �৐�B@ʞ��u���q�c/a�xHRJ�#V�x��I)�	����3�ju���AףnOđ��V���ݳ0� <�C\ּMװNH(�0Q^7�{��.ó��`o�i�D�$��@��/ G�<[���E�?ZZN\b���\Kc�#�tmџ��%	YC�o�}�g��&AW��f4�*�@UtZu�9e[�T��Ȓh3бG5N�N�	�c��'�3w�3d;=DѠ�T��Z^���X)�n�n��o�'Po��OH����6r�9���@���8'%��fcn�4?�c]D��.g�F�e�
/�қI#�����/������3�|ȀZ��0�g�����{��Q��d\{Me/��-�    IDATy����Z��T�[��/��Y��Y�^�*0%SY���rYi��$O�6N!E��jŴ�1|��������n�t�C��ҫc�P9�#wW`��	�x����oƚ5��>\�_gc���p)������Z�|��C�����4�%�Y�����+��CO����&"^�D��&;`'\���h�`�!��߬���G<QD,G��Q�Sz�8r��8�`�6=�R�䳯��;���������nFI�\M��bm���ux���He&	��Ȳꠦ	�0X�RYӒ���𝯝����&��\p~����F<��Gh��*7#`��eNo	}&y�`$�YT��ݏo�E�߅��Y���a��U�� ��1-#��ч���?����1�jj`��%B�Sg��%'l�B����U��ҙ����)���$IHd
H���ʚt� �
�u�5Sn\�́N�ԇ�h�i(p�6����[`� fy��r�v}d�aHϜ]�d�����u��uIn^yc���I��V+I DT��5<�ƶ�?�`���l:�	�?ӕ�|Lz'�p�='Md%Z���P�b� ���P�C��*c��qx�b&\Yy��T�ˊ)��3ב�Re@��.�zc�/��jP�1e�T�ד�&�7G�nI�p[ӊ24����&�,�Z�	�9��ˁˡӱl�)��s��������qD��Sʀe-k�������:
��/4��[/� ,@ӿb�*�R�Fw�?:x�\-	��g��YT��9�q/Z%I$�\�LLYQﴑ�f�����Qb�C�R�j<�t2-fl�ӞW�YruI���̛�^(���.A��JQ�2��z�Š�r�f[f�I?6�X��8�&�CKvZz�ȉ$OԮT�YU�B�=���g�:���I��3ձ���ۉ��Z�ی=��5i4�y��T���S��=��	�uF[�,�wQ��a�K���� ���4V�:U�{���ӴX�x��W����z;���Z	@���?�B��VQ<\e�K������uB�P��ez_U�'����6�L�6m��b JO"�5Y-u	"?;�=��&�4�`;Q�]A�5��}	{�8��c���6�H�)4i��m:#��7`�=O��e�b�hM�A�=��Ri���/_@*���*g�9���U�m�9	4]�
�t�˓�����Ԋ@Þ�[��,ʩ�\�]�mĥVN���b���!#�M���
����OB����3bX�zR��Y�u�Ri�iTСy[���L��n�C��C���]r�E"�va_#���e�<��:����x~�*�7��&8�''�����6	;��r*O\5ЙB���F@Ie� !�ܷ��;��@�U�%���13�}'��U%����!��Y�[ud���_v�ם+���V���_�U���g �U��j���*���b�,\�
L�ē�]��K���.�)ss�^B!�'�0��(?<<<��֩^2ۇ6�h�(��(�j�KĒڮ �؝J�ђ��1�;���hr�~�M�TRb�����6�$nwõ8e��f�`Ts$5k*����/�g��(�XI��8��!�� �H�4�6��	��L��9.f+`j
9�9�MJ���v����P�*.��*�G$�B+��.6S!e�E�+��@��\��ڍR����H8:&�:�g���\ LE*}�lI�V�.[��5�C12����g��Q(Ҧƭ����L���R\v��X?\A.�	G.�׿�)�āFX|����/7c��!�:g:���s��`R�jr�ƘZ�7��V n.�9fǅ=J�7U�������Ilڬ&-����3�?�4l3�S��F��������r�����Iye����>�'|h!fM��à�˲�6��ko�a����0y*B梊�l��/��7?�ͣL�sR)�]Imfa�\B�Q��{�I��7N�>s���vE���*p�Ӥ�V��!?��&�
����ol:Fde�V�V�-)���+�k ���bo��*dPg35���0ix5tڞx�UF���q���^λw���ڪ�mU_c�6T�P���\�nc�T�`�P��Wp�m���E"M�t�6�mx��IYU,��F�=����r!����^G�}3,��C>wk�u1���u@8��D�a �W���}x"�~4h��������T�#Y&P�����p�Q{�/@>d4��Aꬼ���%1J��l�7�W��e����g��ss��7��e��q�����&��#��k���Z.�]���	V�,�u�#��0����t��@߈E��ٓS`*���,.�$#1�	�jM�7��6Q��E`:�O���$]�T���8��F~HȰ�tt�J]z�yP������3M&�V�`ʀ ����GK�ݖ��\���xK�܀�����i��,b	[G6��카Z0���$�4�S9����o�
H4���������50y` �LM�ܱ��h	0%Xd�c����jDO9����T��Ъ��(V/=�U������!�ui�B��tF�C
0�IT��Gm8������7j�����AF�	]����C%SJ��d{x��/E�z�C�T�\cv}���G����i�5f�x��<)���1�'l��}�U0�����J�|r/�����t��y��w��N���s}r��L�sȭT�$;]R�Y2�Lm9�T.�穁k�G�;�L�rmEй�.��q��Ds@gϯ��`����3CUd`N�b�f�&mM�'���;Oǉ����A\{�L���u�[9����m���+������/b��ċ��zxPI#�-p��}����¹1f.�K<�~�6#�G܆5����HQ{Ʋ��u���ʾFgZo��Pu-���25���%�n�ڵ��M�	��o{]�W�#zd(��d��j�k����D����th�XF�}�L��|��.�~�^��K����
��r�x��^���;x��Wd~�;kG�@��g� sjW�ԏ㋷����k�}����GU�8YT@�o5������=��UR�V��c�����ò��[��F�~�P�!����#o@��Ԯު������aW߭������n9IK����3׍RU�lY�R�����I�0��t[h5*���8��{a��a�)Y9��^\�
�����$�S�F�F�Zϰ��%��S¹���~�`?�gɝ_l�J�����&>h�4hW��Ʉ���"�#�U�j�,�� OqW�x.'�϶z��)G���zL	Lkc���AU[�%D<��Z1�J�F�RJ�=�c��F��+��N�!��Ӄ�ߌCnJ�S=��	*�8�4O��\�غM��L;$�ģ�9қ׍TK�3�_`���!��y]S��'A`z4zY1�k�\%0�t��{��7ݍM�u���|�s�DMq����}��6l�<��{�_��L�+��=R�gtt���s��>��_�(K�'�J����]X�n��	L*���E�����o�5��bh�����o���ZU�׎#�I!�K �ja�iY���c�z��!��6��ӯ��g^�W���٫�L>���on����~�!=�t�J�t.&��`K����7Y�m��TL�&b�-G���$g���6���D^gV��M)��:�[٪f���`��}�	��[�f}�� �&*��m�A��٪��n�=�D�e�;�8哋����/�G�@����MR�A`���I�-��9�>�EF*�(׀������!��=H��ĐB�zדDIa<�'Dfc8���ህ3���N�4(��]�ҽH�|�X�uĄ��t�>��$m�t[��M/��w��&�b�'���N�Ъ{(��]����Y_><x���|-J'�ऌ�j�)l������	p�G*���v��ƀ���e�?���Zd��dO&�`����K����н�ɏ�;�iT`JC�m܈+0��.m���Lrd���`ԛ��0�z����T���E���*YS�,��HC?G�1�0-IŔ3��r\LNޛ@�UK����ԙ�q&�uJyK�cj	��rl�<Ef�C�Ԡ$���x>bk�������Z�����@�I�Z�
����W[zNU���b��
��=�<��P��f�<��5L�;{��S���I�>�JY-��%\R��+����H�K	-� IYKt(���:��H��Z��lb�d㙴�H��ѢUs-e��p��2y�t�¶��p=�ν;�m��������L�dO7bx��$\>��ŭ�H�����2W6�:�lQ.��m��h������=t/j��?lޥ_�	�R1��X��Q�������x$�_����p]��.:"�Ti�K� U"���3@��T������\�z]j
��&�i�8��R��$_�\r��A�+�CR�+!Ns�\�y N:�l3%)�"t0�4�VТV)2O��*��7G������������p�d �(Nߊ� S�LP5ų^��b5&��:*D��f�HM}�d����6�O_6lwiC0E��Hr���S^~5�����A��}t!X�I��x�*
�,Uz*"����4k��uddVC��Y�{�`���ݱ�^;b�d �TJ|�y�"C�tV`X!]?������ǞY���&�ı�ȡM��� �,Hh�tģ�Engʺ45��7=�M�`�]W�#C���
��;�m'�ݱ�-���:q6�5]g�u�Dt�;(���j��\�g�p3� +��o�G���:
�h���Ta�ͭ?�GRŤ�����n*;k���u�P�=,U1�l7ʘR���_�(�\8E�4�#�����~>�&��:,�����,�T&��:ۚ�l�a�L�1�����"�
�v�~��(��1#�RHb�=K��T7�!��f���Q�H���G�/���|��h(�M=�\i$SH%��X��	�ּ��=Ɗ=�d�h���\�y���5��GlZhQI5:!���9�G{T���v�g�2��娦(
��[��:VL�H�rZ1�G#b����>L�@�U��|p�X��,#Ҝ@!2�O}p�qڇ�Z�'�N�Gj�n�M�������~l�!�����k��
V1���p�u�c��|��眊���T�I�N��a�o�;�T��#�^� �=�
?��Mش��z��b.�B���	LOŬ�9	45D��[5����bժ	x�:Q WL"�na�mz���~�/��M�Vl�ⶻ�C6��gO�(r6�~���2
f���r�P����~v�b���z�s��ĒH$9:F������m������N�.����:9����#�b��"����<y@�B��:ˉ$�Iɸ4�(Op�(���H���L�܇m���iS'#cߤ���O-+�������O�"	-�NV���ţ��.f����	|�3G�O�<Mq-)b B�VCoo/������ SO;�Z��F���}j�D��u9.C�)�[?��\v�\r�=�D{��T]�z���#%�叽F�n}����'p��)�Y��#�$�lܗ��k��La�x���"���/�H�hD"��\�+oy�F�N	�)�s��赤צQ��I����p�^2T��T�6c���p��_sh���'4.(���W?�i����X���Wq�m�#^�%s����Ai%/:G(A�#}0,{�*��2Y!�(%��!�[�q/2jA��>�d"ʻ�P`Z/i���tR� �N���Y��X��
L�t���b���uj�_�_��.����<w�|��S� %��/�T��R�G��Ƌ9�9:R�)�T�cZ�������ǽU�,�{b+Q�W1�d_�S�I��y��W�))I-+t��M��і�I���0��d�V;�;pTT�Yi�5��rsOZBJl�dH�E4�d�}�14��%iCgL��j?�g�kJ�)?�~K�@�9��¨�u�s���jjd2ZI�t�:�+�rW�7�KF�H�~�����}�K8:0�RMjd�t�=5�ѳ��"�c�d�L�$1rm���}b.A�5�@dП�C
��fI�1Үoҙى��J����B��	]���`n���!����G)���ks5��RrÙ���Ru$%�15�҂�d�L����Tn����و�gB�K�=(?7+6���=t9�:�fyi�0{j���!����b�)d��C#��-����e�.��f��g^���xo�����)�M������$�y�����1��ɯ��)�@��P���s6�����g#F���FY�o�5ȵj��h�7u5	�gF7n��	+�eL0�Z�9߄��1"�k(���W-����6���ѓ�`ם���}�Ⰵ�1w�^�ٵ����́U����Q��%���{�n���$
hEh.�{�����o���x
5[�p�C2��u��k���ڇ������N����E�a�PWX�uk)��K'@�*@�1�V�m&���r&�	Ww�bF$�sK��G�=(@'�N�s�R�U�5n����������[H��3C�Q��P�T��rqG�Y�2{A�a@�lZŔn�%L���{_9��3(N�"U�l���WpÝϠ�C�KS��;%���n�8�H��YFX��W���62^̼����3P���)t��rMz��ۚ3�R�3>3�b�Ri����"�2PM%n�d4ҕ9��4>j2��E�'s�	L�i���~J���"K ��<2*{VNg����6X	SVL� ���r��JcLi�)���n�������<9�$�C��s����Dǫ ڤ+o	'>�<�����I,y�r<˵w>����&(�c��a����}\�)ٍ[�}W\s6m�Q�����t�崃TkML��9^�x|�Ϡ�?�}jJ�2�~?����2�^C1C*V�����:�(0�gެ���~��kʲ�Y��Ȧ���]/~���c��z�ZE3��X�����/�8lo�c���e1��zqԢQ��K�����??�{}�t���TL��Ze�z	��f�?8���eVF��d(=Ac��ŋo�ڵ�����100(2[&v�29*�=]�*�*�[�˗��5�m���dr�=d_��)'b��^1��t#L{��X���dv
z��W��F�iU��q�k���@�E�2���O��N{0�R��{ʥ�ϟ�y�vC��L��ZW�X��k֠)@:�R���jC�֘�N�:��Y3徘HL���yI�i=L�=����D��yu�E:UL��q�7O��Ӑ4 �f�2`i`�dƍ�U�93w�f��Q� <7ޕ�V����F@��~_� *�Z�8��"r��2�^�݂7`��~�/a�y�"wɚ��U0���N��\����s�@96�BoNu2sPyp��7p�O����T��t� � �lNu���n�4CB�U�$)�j�SH�h��H9����h�$.}�H�74Z�ظ��q�)$X�`Z@+��T�3X"����
<�Kx��h�k�����O`��&}�lJ����z��/�h��Q�R�*��?!�6�ϵ50U@Al���~�A�����LR}.*��ql|N0���Py[����2ӕ�Q���N7�U9�uvm�D�4m��{M<�e&)��t��;ǦQ*�,7	V*�I׫��S[M��,�*�	q3��]ʀ#F��6�ꛤ*���^y�4Jji�)ߓZ�|�>�h��hX�&�	GĹ�0����?��L�-������}�P����c�9|ky�#B�%|+7yŚ��K���Ӹ��_�0y�\�J����/ôd�/�����*�[���bh �7����HN�L���O��jH~eɖ�FiB%�QRm0�ˀ)��?�ʮG�jF�A�f�va�M:�E�juJ�Cٽ�|�^pn���
IXU>�=KrS����fq��v��N��2�n}�n���q �wWl3-�{�\G��8=[/}�l�,݈�^Z�Ǟx��Y�J�-2�(MĒ)tbIqڤ�*f��.)n��{�йת�W%���PK���֤���}qUyg�"H� 0N%��:#*_�+M��{��<K_�*�ڳ���@�^�D�Sz    IDAT~�H��v�*�4�`J���7r�n�a��̊�����BI��Il�Jx�͸���ȳ˰a�C��F"�+���������9��<7_:���S�8X黠[�r�a�܊$/��o�c�d�먜��������wc�Dw1SI8�Ku)W��^3H��U?$�R��7���Gx9sSucRS�S��4�	��0Hu����IXq��\�G���B�u��#kE|�T� )�MGySN�V�N�N��{_��k
tPY�[ǻ��w/�e�?�Ӄf7�������s��QL"�RV�I��d�V.�yc@�@m�kk�������9P���g�L�gg�f*���7�J����Ml]"�N��v�}��k�b���O��N�$z�ɤ��s��E��2G� ��K�R�\AetLT�¤R���4b~d=�B���r�i������b�qZ�<:i���eˀ��?'Q�R�9����X1�"�Q�[�'��7O�0���]����TY1p��O��;��D�L=dw|�@��;��˯�6�ۄ���_����!.��)�b�wp.W��n.��u�&�i�lտ[�~��h1F�Z�VJ��ǑI�p���I�t�U~�ӯWp����ڵ5���^�\!�\�����󾄹�
ru��>�/��9j�����k����}��o|x��Ȥ���0���q�KK9�)v�[��jU�+c�x�X��t�ϊ�6y�Mv�������B������Q�EP�l�����j���w���G�ó��6�
8�g�������v���S����n���V����Dz=}���:t��P�W��V�p ����1|�q�ǵ���dk׮��ŋ�����NF6�V �'X�Y�(a�<�M���λ��K���K1^f%�Ô)����'��c�D1���&�����+�E�[@&ׯ��S��.�2@��N��*.8�S8t��H��@��+U���!�J#�ɠ�h�|�_��9���3��Z���c(U��Z�a�x��Sћ�(U�V$��&p�=��+��x-�f;�|�E^w������f�m^��$����~�"M6��0�s�\E��@���]�5��W%��F#�M|Dd�uL����|�噺2���঻���>�j��|���I����2r�R.�ڐ�F�>
�(I�E$+׉ԇ�\"*��H-�#wu\�1�<�Y5c�i�k��e��1��4;�0M�ЎG�d��0�6�ŀ����8��2#V1��*�E��b��W�+�K*���3%�c����L����4�� 0*,�:�j2���$[� ��%:bcoɲ;�|���J0� ���1!���{5�4Ю#��`�7�l*�|6�&�8<����i�(ju����4)}pt��?Y�k�����ڝ�T���x�h�)�B�K��ו�0!�W\t:� _J�&�����Q�Ȥ���Po5E:�D\$o�[�i�,k��EЍ�d�P6���*������Sm�Ui��$u�\W镊��V����r�.�9�E��¨���*gHc���K�:��ᯭw?)���[��K)}3"�'�V�wEֆ`��|h�0�}�
���Fh�K<Ub����3�r������0/�12�J���L�/�AܗU��:�`k���#��؇��V��i�%>�r ��tD|���?��!*㨖�Q/��l�'�����c�>8h��i�f"|_
�ܙ�&8� �^9�%K����.ū�����%T���A'�F4�q����SVФr�k��=�H��2�=��r��G��{j�=_*�T~$Q��4�:K�})�j��K���R�8���G�?�[�S��K�A~Wd�5D;u�SLǱ����<��Θ�� ���GD�]�A�� �����	ĳc�0�ԋ+p���5[PnFЎeЎ�@�e���>i���鋬��O��:�+�t0L����g�����|�R1�
)���\�K�ָX]5�~w���3+�8�8�^��X�"n.�K��g���S2�"*p�~_��R�m�Q�;���g��5X�M��ϑd�\���~~���Dr-?ܯT5PMGe[H8��*a�@?���8x��(�xg���k^��w=�f�V�i�'��#Tt*���>n�=�5��l6C2gH��U��8T�A��j�j�pg�|j{�Jp)�u0K�fk��:yd�o=��B����1�"�J�/�*�u�~T�8�>�e4Jt3nI<��x�@��h��J�U�1dŔ���F�ŕW��=�6n��y��]���j�)]}�b�v�����y��9����3p��ʔU�h�j�:�2w @�#s��G�P`�ُ`��/0��O��{�p��|*��[����q�1��r�=/�ˮ���[���A\��`�m{��]�B��B,o�$��a`���|/�)#u�[_�%�;���p��@6UǑ���y�8Y�)��c���s��v]�hN^:E!�Ǝ3s������ff%q9o�`xd���& ����+o��^��O;��;�f�l
o���]r�{e5��X�'��4�V�cK����i���=�I�t�m�����:�KYxe�&ߎ׋�a�6EL�n�\�}<�;�y����y�i��WOǞ�o�3͕������#ƪ�S�Q�@��#@�1�&�M^su�V��r�2���������r��͛6c��:�ªaJ(��Ag��F�D+�j��|~w�Ux��$i�)��3?�SO>=ʼ���M_�eW��6g���R���фVx����f�V�D?<�,�w[p%�g[�<�\�R�[1_���x�ie��4%�\���nw�-U���K��G���W_���[0s�T|�s�����0�����u\t��*ǥ���wzz��)m70�a5Jë��`�}�8p�t��V�*aX�b%����cd�$ILOO��}r�&�I���atdL>�T���W��j��m�����c����I�c����쥾��p�-ϣ�C����cد�i�� ��C������$G�:.řv��܌tьSʛ�>SJy	,ɤ�8�#�E�6ʛ�QG"��r���2�$����6'-��Hj��r��qx�Jy�*��9��@��m< ��@��4��0�W�*����x����V��$�RՐl<��wjk�##c�u�2���H��G����x��9vK@�a�'sx��*��>�#���硿 $��W	�P)�#uL�*�z�Ȉ���+Z��=�N��|�:,Y����5�`%�D�.��:Ï=Rr/��f��o�6���vS1g����չ:�^y�ʍ�����1�<O���q�L�L�F��+xm�f��RF�C:��V2��(�nl�lvK��jF�K�@5wty�`KgZ�p��W,	Ti���DͳXL�4)u���Ull�e,�뷔5� �&aM��)v��������2]3uJh���8C&���Z1f(k?��N��X[���}O2B&�X���#���d_�l�ӤΞ�"E��Z���C�/n�������5퀼yU�n�~�)�"g��r�b�k����2G�#*���f���Ht��%�{��8�#�ߞ�`pRRA��e?�4�.T�y6�(9﵁��eX��J���m��|5V�ی��H����<O/��U=����%�$n�`�8$#1d�+����9j�/�I/��S��s\"��KZ,pFL$�I�Q5Q��fKr~N*-��QتKU�����I��f{��	����=�O�Hƾ]i��su]��=�����2n=�]�&���
���*n��H�XYuf	F\ңRu�f1"���"�G�݃:{���$P)rpd�TƌpQI��4�:��I5[+��<���̕���/΂v}�:���7�����F��bL�ʢ��,Rߊ�$`���I��CJ�@�6�~��=�~mʃ��$9�L�.���۶�i�;�����>�r�}�W������~_�v�� (%a�ji�YG��a̙ǅ��$�e� S>#���������^D��E�s��w�Ɔ��Uga�?�!���UB/�$�Z0U��EuV5�*�bJ�U��Y^��(�V)���P[�ĬД*������t��-�9���ƥZ S�b@�����L
0�#�W��h�&?+	l�)�u����2{��9�)a5S�Ӛ�tJ|�fЈwŗC�$#��y��*sLK��݈f͓jiJ��T<((�<ψ�h���ٞ��%*1Vr�ڈ�j�5�Q��Cw�Y��(&'�������[ŭ�=��z�d���z��PLhU��{��w���m����?;f�T��g�=�`�D���V�$�=�T��G�]��a��݋{�P.�)0M�q�a���o~3�����e��y�Ɔ�- �GJ�+$��հ��~��c���j�����YDeDm�|�E|�ďczOLL6T��?����2�B.���MI�L�Z�҄�����O���K��]Q��zp��g�%H��7z�@�$�����q����ŗ_��g�k_>;͙$������r�+��ע��� W��bq��ۖ��-��H�gLE#u�C��6���~^4[g��Q�� U�m�� 音>5��o���k�/{)�u�\g~�38��cQ��3gZA�/7-�����V�t��')�%Q&HZ{"��$����g������ס%k<'J%�y$�r�g��wk뤑�[����	,��\y�X��2��_<���W����Q�ƛ����}��4�׊�w� z�������G6��ئ��������{��o��^{S�)+�d٧M���������q�T�U�&*��9����	,_�
���+V����f�k�C���~{�g?�O��2ro�O~}7�[�b�����!�ۇT!'2eqГ�1�x�,���$ Y�m*0���"^�#֓�Ö����P��IE���Be˨ S���7��z˦�I��Є�U�(� ��&孏�	0嘔���F
Y1Ob?��+�Ra�L��bڭ�|)���6H_�1�L �y��STޥ@đI�YO.t��aANL�|�Ss����u.�26F�h�E oO` [�O��2��5+��n�3�
'V�U%M�K�)G2��������^��^Z�H� UN���T�+ÿ[m�@'�5���r�Q�{�I��,�18�Ɯɷ�|?g���&cN1\�{r#.��lm ��IՔ3#Y-u��R�U�˱��R-��Ry��Z���A��r~uB���=s�˅O��A&����`��ONX%G�˘	�E�p���a�{V���T׏i�}����_�������:�Ѥ�~?�U�]�3��8�=c6�f��ߪ"��"o�\�@��A+��*g��M��rVX�Ku����[G\ʪ��T,�ɨD��"9��/SbIO��d�u��Χ�
� 	l���ū��U�Ѯ��Qقb��=v������������*�dUH<�J��P��B@(ՀMCM��|V�ڀ���Κ�xg���7�l�?�����ӨVPI��<��é#*H2*}�QJf�q�Ȏ�@i�6�Uǹ�H
93Kek��#J���hs6r�h=��2�ܓ���m��`�1g����Y���&;9b��y�}Jv�Ɓ�o��󯼅�~�+hŲ�&���K��D�������m���X׊�58u:�8bJ��}٪�K�
��@h��h�=Y1�yײ�hi�7�D_1+d�X��r���HKk@�p�i��S��Ą`-�
~��3�e\_õ������2pu#��K���*���֊�'k,4{տ�.G�+�?�U�۽L]�0�������I��۟��;�ZŔ�Q�v����Y���+hF�2M�$'��x1��F8��QM�*+5��*�̏�UW��{��`;7��@� ��Xݨ�/�7�-~�`�ӹ+��3�e��*9����@�dIJ�}�cIx�>s���)��m�3���Ҝ��E��
���9����2�#�2�E��M��M'��H�*�K�BR!A:E�*�J�k7��t� ʶ.��I�0�XGb��.s-;�k�R^mc����*b�8
���M��$��G��)���*���n��	�m�1<a�^��g?��%��~s��X�v����?��əȊ˨U}��1�[3��ÕB����hF�Q��Ԓ	\zŝxe�z�]��d�SM�h�=�$L�L��E<�tg��l��;���;�4��q̜��:.�*.}"��ċ�,h��t5�n��=[6���eU������5��-d0��������������L�ו�;�1���g@�C6������Q��a��:nZ�(z�q��|�k�c�Y��J9JLL����u��/��X����L{{�e�rA:�rv)Mo(���(�A.Q�O��
�:d��R0�����P��- �U[B��'��?�k��W�NFp�O�)�:=y��*G��ox���z�5)���O�8��'1[b0� �Hy3�q��٧���1�#c�l�J��\����~�}���2��$5�!�Q0��p���ફ����O���=�z�B0�a����_�06�G�h��;i �}}Ȥ����1�iJCk��`���8`���gx��j����1���	^6�J�mϐ|�.�H�-����{���Ï����wWJ�n��|Y�/R,�0�����w/E$3��~dz���[/� �2:O)mf�9�&+�]�"��tФ���C�7�v��λ2�Ĺ�܌SJs�&�[FQ��ǘ��B�T�JP1ɍ�J��(*�í�20e�E"�Cjp"VL)c2c�ZW]�̊���f���d�Ԫ�\	�c��$Y���oI�s�B��k��&�Q�[%$���)!H��7�����EC��Ht&05_�/p&���=���(���W�x�R4�1)G��/���}��$���]���8 J
%�2�u:��tpұq���`�����P_��������o"�� /������֪q�"{z���{b�t�0�v1�9D�%{��Q�v���+�c�]�%t�
�=`�1"���_.�	I��l�V�Bc�UI\�uD@P!�s�3J;�|�m/�~+�/:.�c��I�y�3S,Θ�ޥn"o�����߮br����?v�ދ���xgy�lfGE��v��Y�rQ��<]��p���_> 7٢#��?����u^	�����%�>qj*�I�D��Uӓ�n��0��(ڵ1$#5�8{
��c.>z�a�?w��;q��)pl��7�=H��l�7�RX���W�X���X�+�b�!L���ت�5e�o4�2�m�����j�����ڠb�$��&k_:����s"�c�CM&(�cG�?��{{��={:�̞�9�L��m�`���Lʢ�@u��y-�2ٺH�5��߼�U`��a<��+x�巰r퐀�H��H*�NL���t�{ Ğ�4{��:� `��Z^��*{�zf�����p�/}�u��&#���G�.g16���b�����A���`媇����?��'�-�E��sX�A�њT^��@���*���82�d�v���#O���E� S��_�I���ʽ�#�����A�$\���4����]o�����FL�y60��:4�C�aZ
�u2�ݹt�����a����p��K�E�%3�X博^��ۂL(�R:�Q��3hr$]�Iwu���9����npJ��Q~��-��jg�;g��?%��=�L��Hyi�H`�|���<+ ��Ođ�D��*$�H�wD��l�>��O��>1	�r�M&��Z����j(Τ��H��7Ly���Y�.q�)��xH�����Lu$��O����;���L�p'0mUk�P�>v�VL���)�;/�����S�6;(d"8�=p�g?.=�nw<����UX�jj��o�6����b����:�f�>�T���<�Fs�U��oxw����0�f�Lh�D���:d�9�D�`�R��^-����[貙C,�D2E���rm|�#��� �D����J��^zs�.ys�w����T�z�2�pۣ�U�C��E"�F�]�    IDAT�����SS���t���n�TT��Y�1��*���b�����/����wq�]O`��`�ys��3N��ii�R��;\�����c���yl����L��K�|��o�Z�@,�!�G>Y��x&�w 	&����I��п\� �S�?��W���O49��/.�o�D.�W��I��ћS)/�n�t�˸�ƇPk�K�b�ME������VL�n �:��qq�^��v!`���5J�i�#�u��F妙���o��l5�;��xᅗ�Ϟ���5��un/=Ni~t�C+𧛟Ć�(ꭨ̌��UK(�lDmlv���}�4,ء�}�LG��?
 `�U�&v��>ee������57܌�W�;l������o�]A΄��cm���X�����"�ӃlO��s�б�#3��Uζ�F~�PJ����iT[����=yD{r�'��"(�^���(�+ouh�1ν�NoyJy���xݦ���W,`J)o����C�Z1m��&�5`J)�4��*Q1�]Ć=�h�	��=g��lEH��������c��u�9�$}��6��3\�� �tJRl�O�7�Q�����!�Ռ.�T�7��(#��c� p�_Ƽ�aS�@�b�U�]o�}~�����&�0{�&<��=��\�wD�=*ǌ��%U�IjL��=�&�#������� ށ��|�L\��yc[���
����8����k[�D^��$�9�V��n���XNΪX�� �T�����Aw����[�� 1@ο˧��HN�ڤɘ�e��5S��*FT2�5Xt-A���F7�7HL-� 戆�|KK�sE�ʟ�Xjl�O���T�� �*�S[V�}pߓqBtU��gV���уv�Y_8�3�+#e�G_�7?��Fڈd�Ir ;�[XRWY$�[_1��c���5�T^����w���\�1W����sS,��C�!N��:�y2_�C�aM<!��J���61kJ��cg|򄣰缙�1|Z�(I�=�����N-��~7� �J�ѱ&F���_]k��n�&,g�z{5�^�[F&�n3��g�an�FI�M�/wv0ݯ���RCN�L7�"��a�@/�M����~�L�:e S�1e��=1Q�q�0��|%�gfy�VH���H]#�	�GJ�3/���O���o�Ɩ�:����ؓ�>�dZ*�bc}�r^وV�M��Gv�׷�E�eo�4�W쀦�%a����P�QRN%�2oT̐��i�TC�6�B��O|h!���C1�_��9��W'p�wa�6Z�"��Y���J�GK�g��3��yZ����\oe�E=���1E���A��¿���e�;���}G<Ĭm(������Td���lc��c��v���0-�����C/r�v�!��p�o�ݏ��F7�/"4��x��Hb ڬ����F^���1tSt"t�O������3E]"A,t^Fq���00�B�U��Ka��f�2�Ѡ��r`*-�L]Ŕ
/� ���4	Nk(�w��LY1ph��Y��4C.��^��ظ8���i�X���r��[���!�l<�"G	��1�v#ڍ����9!�m�6V�h��x�Hx9O��]	0��R�o���ᄃw��?�R^��f[��̏���ﯾw?���6zsq��8����-�`��/~w%V�ͦ�*{�s��N��"1t�*D�A�Ge���EǾ��coB����S����oê�ԛ��$%�eS��6��E��[_:��Ak����q����+Zi�a�|�GaL`r��}�o�#틝���4e2� �k6�;�ҷ�����>�8{�T�|�M���JT+L��((�U��)_�Q�H�i���/�����}�&�6CP6
7����]�sY�)n��	�씣j��3�8�^�/����\���z�?�4��cg|�Ӱ��"'"���܍���W���R1M�0i`:����Kp�}s�)�B(�f�z�9����?��?�Ｂ�Tr����|O%�>
ә;�OIP5!�|q�\�_��w�!��_9�9�(fL�H��oX"�F;�x2���>�?��-���g��j��d���9���v�7���ġJ��[��
�����!�j_j�,~�\�W|��q����'�dG��c��GW�/�>��z�f��>L�LiuG��K�P������g�9s�I��,���E���镻j�W��̕��� �~�<��s��;��׃���Y�͠0g�N�
���Ý��Q��G��μ9��G3%&ج�r�)��.�(����t�FdTL�'��Hy�h	��s\L��R`:Z���@��4�Mi�=�C�Fy�.J\"b~T�(���Z�g3
L�|o��x�k�� SVL#Q�cJ)osx�
G�х�e7�NhWHo��X�	��6+M���H�N]H !�82�Z5gb����p�jD��]@���EC��"��HYdJ��6��U0���Ͼv���C4'P����:�kg��8躖�S����I����݅�_\�H�(I!��E�lR(>k���s�4���q�q����B�h):�
�W�\OvW��=-��@�u�mD#xg���Ͽ:���ǑY�� uv�
�J�u;H�a24��"+r2n��"��J^|��qm��g'�)ֻ�J)װ��\����Β1���7'�cϞ�%�U���?;y�VVx��1�J��ez�]�[{m5�w�S�쁙�/�5-�mh��%������%��(�J������#�E��g�4'���KK�v�cx��-����uT��H(�SףK�,7ٺk!���D�@�|0���3T�@���H�.�w���#L��=�4;a��C�a1��į�^A�<��7�T��E퍣?p������!��(�6�]-���5W��g[�N��5��{.�+����5k6b��-�^�I��q׷,g��%	������z		�7�c�Rqd2IL����郘�_���<�,��s�Q��蕾]������e �+��g��R�#Ml�<��W��}>�7�ل�Z�V�l"	��I#W�b�v�2��g"�`|��K�������� �;_d���[2�u�./�2��ϑJt*��f�m�:!gz
��K�#��3���qԝpmI҇����n�u�#=2B0�J������g�[���E$/��n�<�g�>�J��[�lN&3@rَ��: ��{��~+����o
��T�=(�˝���Kw�oL�9S����d�������iF?��)�k�^�͕�ӵG��wqzn%��^t�Y�cI48#��D<�@O��A{���(U;x��U���'���~7���=w�+�:�������R�ٿ[� �H���nM:JF	P�S��`�Sh/~2�D֤�$�9Š��'�Qj� �4�+��+��1�$b~D�CTBN��5����������3������� 0eŕӎ�!��M�D�@&C���e��݀��V`Z(���0�I�AL(4�rF�r_D�����V��YЮ#�.���qw��_8�I���W���v�^s/�y�yT��1�p����g�G��� ӵ����[o�G��!����ù�<��<UG3�N7L��	o�o&c�<��|�Kߚ��t�|y-ƫ19��IvY���6PL�p���/�i�Lu&��Y���c��N!�M��׃g�5k��]}�v�~��Nn�e��{k7`��5�7�&:�y�98��#���������k���K�bd�!��QO+�d�	���qt�C���R1]`�T�y�7���+K��%KШ�Q(�DI�rV*e����&��ɂ�>c��4}3Љ���ꍸ��G���/b͚5�����9�g� �Y���ҍ�'����^#N�ž��6}��Yp����+�t�-��۩��P`z񯿇�w-ho,��6�~�y�\�
�b�lF�����,�(R����U��8qfr�PΚ�!���އ_�/{��F���q��Nũ�:E2�n�U��q�͏�����q)R-(Q�C�f�$R�4�~���}`*y��UՄ_�}K6E��$d��u��C�s~�ٷ�����/���AoN��87s�������o�a����r=���d"���Ƈ֡6�����³?��f���J�T=�(H1��(!�ǒI����'LW,"��%��ƕ7�!��_����i�A��gn ��������a��T����� y� T��P�(0e��7�!H� <�����H�d�ǔR�N<&��MG�#H�H�~J��C�θ��r��ͤ�Ǵi�ׯ�=LAŔR����1҉f�HN�Պi�=j��E½���DG���4�)	0�T����;򅀩!�]�/k5h�0���WFě�@1���O�.sf�7�F.���`���C�����x���X���Z'$��&d�pcb$݌m�A�!��6�-����b��b�*�'Aޮ��&{��S����5�����<4Z����x�⟯�B��d���� E�ZL���(�b�U�,a��'��}w�.;�¶3����*8�41y��GG)Cϵ�}����"z�)g|�x�����"[(��Xq�!+G K3��%��Jh�f���^�/�L���Xg��@��GK�D+�40j�Kg�����P���Ӻ?�4�����gZa}�b�a�.��F�@A���00�?��Es��$JxhD������xI����u[�Ć\w����8�ЙBPsO2)b>��������1���k�gьd��e�7g�%Wue�+���� �0 ���	6�̀1���<�=D'�	6�$��@"� �rh���Օ�{U�s�}U�������:U�w߽g����G��l-���G�D��?�ј����씍�a�cA��
Z[����e���7*R���Kt��Z��*�?���Aj�4,Mψ���	�8h���g������ �@m�Ca�[5����s
�q3ڥ ��u��ƚ���T�����2K� U�q8_�lq&7\f��]�Z��5l����\ܙ���z�\6l����V���k�������l�"�e뎱:R�Ț&��k�?j���n�1�^�u�4 ڏE{��L�qbVЧwC9�R3Fvf�A�r�!���Td=�8(��5�=)���2��'��)�y��E˨�p�m/�ɗ?C��?���u~Ua��� ���㲲�z�Em��-��e��WE�\w�h���*;d6WƘZ�k�ڔIFqAF�2ඉd�]��b�s:Cn�;�g�f���f��έ��[D��3�G�k�þ���2�Z2�]��7>���� '�	G,,���l�>Y�Ӝ^\~�I�fP�FW����}=���@(��:����yP�s$�[%(��73�-�5mrx���6%=E�}�V�����]��1,��t�[L}ဌ.q�V �D��@�$9��R�[P)/gLYw�N�����	4���*x̞	+0�CF1�U�JE� �j�)4��1e�*�'I#E�}0����0��8����®�	
$t�e��S!c��$0�v�8LC�!cz�l|����{�tG�����%���4���qƑ����N)o�	,\�7��|�٠0�P��|����諧bboX6m{�HGL:R���nۦnn2ݫ�����������Ko��$QqBE�F�d>�H��8�����8}��]s.�w���7c�A�!���RZ>^-�@��-�"�
]�8G�D0�bLr�U�}|����c�9I ~V��-���G��l@f�1�L�i>C`�wF������}s$.�k_1�$������ʕ��ۮ8���1vl?B᠀g[ �n؊���D��&10T��O6�Օ�0��Ȃ;��_��c�jhDW�f /�܎�����:z&a��I2�F�/n��|Q�AFG��eG���h�FН��[~��vK	��)�/�w�ށ��+ƌ�G*�Y�Z��I�8�Nց��3F�T�c�b��	�7o��	��J�*���<�s
�j�&�]����?�
��N��H$	еi)�n8T_/�hVnd��߻ G4S����a�T*x���G1e�x�*ed3#��ܘ̧%;�!�HI�+����U`�5��p�M���G��.:�IF�k����O-Y��^��0�͐��'��á�ں�� �N��/pf���0ϋ���=b[RMyd��� ��%׶�lS���A�6߹�+�=e�t����ԁ�q��x���阈IS�"IY��dt���J��b����Cjf7D6��|V����I%��d%�a �l��W��1-gZ`�X.� �����b��2�H�/�iyG�"��@ E���tuL�H0�cfh9ofL���p�r>�AH�9ch*5��j��e��@3�����i��C��}�.:�Dy�^��G���:���[s������/��G^�����v��t)���Sؼ*�^�"�Ŕ���e�;�COXe�[�{k�̲��;������\�A��P�Y��P<� 㪂AĢQD�Kk���Q��N���z�j�zQ�w*C�Q��)cq���'�H�wYc�>Z���� ��4�Ξ�g�� ����ށe+6��u����Ṟ QsKeL�=4*���:�r�M�7�f�t&��G��g<�0���Vɟ�)(�m�e���H#�csN>���f�H�0!V�i�>�vFɞ��AÈ�;-�Ҕ�mN�T1HǔI�%U�Qe����l�Y�F� Ϊ4�R)��k�u�2;m��G����O�i!�upߑ��Ǜ���yϾ�!r���n��1�"d2T.�l��C9�����m�#��̧[�����e�M�e�y�4�'�J+�5��V�gTb�$�f^�Ո�t���^���;��}�I�c�|�>�}�$$9i�lq�0��2�LS�5	ֺ��qo���L^��?�d_i��tmz���m�'��Q���Z�,�k�	�a��W���a��\�(�j��x��O���ٺ�kܿYs������ơ*�s�&+�b�ٸPc���H��j�2zYo-�}yr�ܽ���� R@gG�y��j�U1+��GѬg�����q��cE����MN�Q�l����?��W�BiY��ą��^W���+',����i���6��T�m��<2f�jݴ֚S��ǚ�>v�wbo!h����q�HA�� �
��=�6��l+qu�"��[D��3'�p����}��7y󔓲�������6�^a�y�������y'����rt�������w|>\[@(�'���)��ݘ�S���ޣ�����Z-���,
��3�
1�Б�j�CSZ_�QC&.E8U�5�̋�7���jد� Ǧt��D:A��G�ʲkGrL9cJG]��(0զi�Y��� R����t��vU֠�2�>��y2�| ��O���&�AaLYoeS�K���$���Oe�z��b��i���|�րu�u�H7�8���{�4�l69�����ƳK^K�T؇3�����)b~�����A����b��a�\�� ��Mq�\\���e.S���k�4A;_�M�����?��1>^����z���%'
��k畚l-|s�2N;f?\y����Py}�^~7��^�d��~�!��\�[-a��uh�ʲ	5E�N�5���H}h�^��;��s�k.B"��{�p�}����Uh���@I��/�J	���8`:~����"����k�^����<���7�_�*&L�,Q	��z ����$_��?Ŋw>��^çk�cG��?*�:�~�$����	}��,�(6�X��n�χ��&����i�#ҀR��f|fG��t�4��K;���`�Y	����<� ������x�M�$�t�Z���LV2X�b)��(�P�������W�xc�,}m�XW�C\y�ٸ�+���2｀<Lx���"�N������$���z���ˌ5�� 0=|�1%;Ç���Nɲ;�C��m� 2����d*%���O@*�%͏tg�4��ڈRx���-�×N;W]v:��B��ӗ����_�p1"��q1S'O�tl�K�    IDAThp ��~���f�;���'��쉜�����2�lx���ΰjŭ{��Ij�l	�G/�c�r���c������3i`��������L��1�0q2����9X�X,#3��?�4�=P�Kۥ��Q�1��
eL�0���Ϝ��x����VsQ����)j~DƔ�T\yM��W�`J)o��i�Hy�k����;�����'.���ϟK�6�Z����C\y��j$��{�����BX5{�t��'���rv3�S.>��8�����B~��AmO�ui�G<3{��&~������MM$B,��2QU2�E��YL��_�ݧ��S�>񣇀�$[��j��_��;���'(W|��*�;�������C�*�gL�M✱+��=]�6e::��:�	7����0�lވJ���d�&�����;���69��*�p�*,\�B�c�̘��N?�]���Y�[�ގW^ۨ�t�8��z���e�,/��˚,Q�pj�Ŕ��S��l�d�h=a��^ceC#!�Z��3��)������!s��#)��̀1���5!�����̵�E�ܘ�,ִ��dIF'��6{׬sy�m�u����d���r�W��"n��i%�X)��Oτ�]���.Ƥ4���⠪�E�� ���b<��-d�1����$�n:g�š۸Q[��Q��S���t	5Y������X:�>�
Bt�T#�ֽ�������Z���?�&�Vz0�P-��gSԭ�Y-H�ՙb��8�x�8`�=���H�*�kC��ʪ�ֆNZ��<s�G��PyM�I�`�{�[ o_h�v�z@ְr��n_۶��.?�*�������l�K���e+Wap��|Ɂ/C ��IfeT�rV�	��H�I\��g2����qb ��,t�_�<z���Z{({����b��W-c�g�f�ڙp��t,� Y�u��2�E:6�"�,�#��}��_.<��N#!�(F�*L�_=1��W6��`[>��F(��r���*�c��Dk�� [S�Z�}���.55�-��9m��-��������i\�k��l#���D��/2�?�D�g�^#=�X�׵&u�(�aքn���gZJ�m��	Y~|���r=��jlp�p��b�]:�o�:�N��1�����t�0pՏ���VmG 6���4o� yEwR��s�A��#�w4�N[#Цx��k �S"���AS��ڛ�a�6�4aŅRlSΘ�1�)�:�_2O/��"\o�����S��ƟAW�dR\yku�%vQܬ�pb��q�dQ�H(*F�QL���I`ꝇ��1�4D*D=�Cv@͏�(�p��ʘC��J�c�f�Zl�2G'��O�í�_ϡy��Q�k=����_��l��[�y/,}Sr�:b��sR���`�v����a�
�����H�Q+!��C��W�8��2����z[1Mf��<�y��d�X��J<�«X��vTq��le�H\%$��b�I-��Hg7W^tz�հ�%��pՏ�����B!���4*����u$i7�
��ض�C!�䲃G�껗��#�V��0��w<��W|&�1*�C����Ā3���M�U���Y�����l%�.>�h��{̛7����zhMc�#&?Nk7n���ǓϿ�W��;F���#�H&p����+.F���͡������A�E4ُt�S��l8uW"82���(s�5�hֆ1y����Z̙2��n�k�m��>���G2�FK��A�qfg�l �\G%��"p�c�ර��7p�%g�¯������<����x�e�cOtIc���m�(hID��5�h��T�k�ǡ�N`Jc!n��l�>��N���O��Q�H�2���G�x�R��"�c���qT~����x�a!.>�|�ʯ�+I�C�0��K��?�]���D�FG�$�(��Q,d�}�ZF6c�=��Wx�Tl*�F���q���9��S��C��3����`OȿE�	�h a�b��՟�ǃ�=��L�[����1C�G|n�F������߇�Ƅ���ӌ,�R��b��u5���-���Jg}���q՝�cS�2�A3��+���fr(���QR���1u�Z\{�c"�;�4?���aL��1�q� @ �rb��<$�~��8.���Bq'`��W�;���Y.3b e��{K�V@)�_=�|��/��]\���s�F4�̲���H���?>����p$o��`8(�D�����Hy'u9����i)Q^�lEa�$ լ;T�|������p� �2� ʕ:�F2(���VA�����U�b�ЕNb��]�������@ �}rÆ��^���p���`��>y���f�mqSw{�%ao�̘���<�i���{��Q��߻/����=c' �ݣ��2gj!'���լ�i͛l�h0̦�E�o{���Z�S���jQe9Ր�U��п�8Ơİ2Kc�l�5�S!��|�6t��46�[֌�b��k���Tq�6L�-0��y��W�tk�d
)�=y�'ѳ�����!�Z�^PD�4�W]r�=~w�6��Dv.N��p]ozj�{t)�����4)�9�(&�A@��!�I]A�n��u�a(�u7��j`݂R;�qg���kG� ��ZWl�S-b�=�o"��H�#C�V�V�2�6�ו'�93�b��q�߃��N��됹T�@mu��x��,�qm{̺���O�{P��ֶ���bD�H��u}�ZM�#��6�}�}�R�lC#9��a�����>]?��R?��4���Oj<�$�8C�$��_2�4|����Z�$-h��`P>�]��:tO7r_+ӗUcA�l��+�=���蹠�J�/G�(�-fᔆ$z����g�I�0f�z��1X%�t_�j����xM�p*�� ��nR.ʸ��؆��Y�#6��KJ��5@�m�hW����M��3� ]��v�?�(s=�� �(�4�<v����f�mc�vD� N묮2��Y��Fs���a�I)����ה�1?r� �L����յh�zP��d�?b�Q���ŏ��$�KT�)-��8��5\���p�: ܏Dw�0�������.�"�<���Z]�?�mi#S�;+k7M;���GX�6��e5CR��5w�0�/]y[����|/�~�#C�ޔ��z��q!Cz�(�$|�*>Gs�i],��AeL��� ��pF����z��2�0��� (054	��t��P�!�u� Sf��:;e>����W������Tb|���5P�;eL	L��Kƴ�t3��	L��)��_:z\|Ή�\�r~~�=ؼ��|������;�����v�Ѕ#����.����0[E�4�]:�}�f;.yO/X�R=1Tv���� e.'��^���"�<�@\q�	���h�;9q��è5�D9��S�{"���Gc�i���]ģ�8��\g�FF��Z��j��P؇iSƣ#������E��o���?چ�/,��h,.[�2(o-����3�����>3{�C�t�6o�(L��Y��{�쑐�v�L��m5lپo�^��?�X\b7m�"�DG"���:�~�L���0�NRӇ'�l��n��Z\\y������,��Eh���cW�\D(�D���.���/�-�sb~$N �C���[��!�s.���a)�Ŷ��Dw��-7�G�{���P�5E�tم��3�F�C��<����o�[��X��D,�%C�Qp�ӽ��ّ{D`�9��hU�b�o��Jd��5����{�5ӧM�Wl�qd��֤��YDo�oo�/.}R!6E|�d��/�����tĂ��L?��S���(�ȗ�b2��'P.�݆Jn {����o���LwTgf��˖.��iS��Յ�ӦɃ�n��˥���f��@��@�PC�|���w>��o����L���`�9ӥ+ɍ1� n�w�yt%���	��E%څ�V�zC��[�!�ڜe�KO���\C\�䈔7�0�b��P7m�����9�!�)�2�c�j]�-����'�c�\/-���V�A&0��)�����F��J�N���#�{�r�TX2��E4
:cJ)/ߗ׋�E�q�	�7ֈB����`H�������]�Xbլ/��J�5�E��\0�7ݜy���x��7Pi�xg�|@���'�P3�I].n�ɕ�35aL�Z�>9�@^�8"�����L�RM�����T�!��jL�HG^�ё�4�v�c�H�O򚏎���H�m��Ɉ�(���ʝt�j�G�x���w�>c�t�?�7�� ?�!\��;�x�:�с�����"0�,��{Yi�ȵ�Ο�$�_
5�'`�>����U�y��2zBJ)(��� �R\"ٴvO�f�vm S@�u�5�mL�c�v��Y��ۨLq䝞���|i�E)�1<����G�.��تv�2��v\L,E;�\���^jy�����8��=NF{8�%Z�#C�o�~��|k���WC8�5h�d�5��Yܖ1��7cJeF/� O��rf�g(TRǢ��3���`-@M����WJcXמ��d�i�!¢�*��u4jE�K9����Ҙ2q<f�2����+����u�#G*A$��_��c��@��l;����_Z��(��ԽFYo�2��ګ�re�ۆ2�>���"������wF�8�0*�OfG]aDy&3���M=�*c�Te�!�y`f"�7��u��]<A	����*��"�#�u�T�g�w1�g1��e�M]f��)��Rv��L���/�S�= S�}:�%���:��f?������^�����EbҀљR6��{¿�\M�V�$�D\ymڀ��%��Ua�ok�A]�x�ƹٽN����kȥ��vf�[�3�mω9�<����-��g�_�휦�
v\�TPA�0�Y���_`��g���d������OJ�����1�2|�������X���q��d|^~ͭxm� ���w��G/2�����L�'��Ҥ�&�`���h"si�ԕ��eHm�T���I���A� � Mb����1���z\����	���"�H���b4�'��*0%c�g����2ey*`Zaf<S��Ad�!�5�"��Ѩ�����:2�K�iG0�Z&��� �Ŋ �DW�S���j��
�Uk$�kPY`Q˱QAS�z	!�5�8� ���_S��_ߧ����#��_��}� S:V�����ց�����t����9p�y����A<Tǔ��8氃pȁ�c�����_u��j���dp��O7a�a��A��	4�ˠ_P:q\I���V�{�I_�e��nNR������ǿA�D��Pێ�$Rq?���k���I�����5e�p/\��8��"W�ޚ� �w>��?,��h,?A�HG3Ac�2zce�����/L��.`�l�,���Dܮ�15k�c���0��:ʵ:���3<�p9>Y����|R���>�h\�/g�+�rC�a�#�|��o{��U7�p����Vf#��jU@���b\O���;���,�A��UĲ��q�� �)��C���H�����x�u���;0<ZAG2��:_?����6}�r�o�᧖�R�"��B��z�D���ܛ��?��f=�:���,|a�I�*�����z�u����+g��+dK��U7-���������<�-CYl�I�s2�w.���w�aaQ�K&��~�;��2JN�R�xa�s��3J�Q�
�{vn��;��cd��e5�ګ˱u�&q����H$�ҝ�E��L��:ՍfKxe�x���ؑ-#S�a�H�J�H�Ν�[��3&�x����;^Ľ��7؃��^Y,�9dg���t��hN����5r|���a�1�!��4�bc�F,d�d��������.`vpX����U�4L�K`�s���c���ʘ�X�� �{:`TM�/�������$�r����� S�k��9����ˤ��u�MRꃦty�	��8�a\���o�c��0[�X��;X�a+�m�!(���)�p�|̜>�J�M��E��?.B����לs��r^��L'w7p�O���&Ǆ���>3R��"\"�����d"&���'���5FS�f
:��k�V�aݺ�B�>k���sV�S�5�����L�"���1^96�^�h�=�Xf��}�q`LZ�o���&L-[�߅�������)��l�B$�r���(�2␘qv����T���͂]]��XY��d�\Z�pY����J[��6[�X�Ԙ�g�����r��>G��}��rj{�	�{o
L)r�z��̛)k�X0���ڥ���֕��D!85��e��6)�o�{<�x�.R��Q�u0�M<zQd���l�m�>�϶��w!����$ɽ�L�d�*(�٧6ONS���j6�OS�{k�ۣZg�Eh-0�#F��ϲ��v�\<���6X����r�̐IU��ZC��Be��н�8U��"��c(R<�t2��T��;��'M��~��v��?�����ۚ���1����4k�5"�熚'���0�u`4[���۰v��۰7mŰ��jV����@D��Lp}���M����'��K^u�բ��[�<k�e��ހ%Y+f��_;5hLSŞ�;hж0V6�4� ��=鰂��F'�h�F0���U-�Fy3'�qѹ�����$Ö{-�+��4�^|0j�I�~x!�m/��H $��a���k��qs����;�9���	B^h3E�9����j��GRY�;�'$��Y�������S�.?ߜ�޵2l�J���c:%Ҥ��o��^*�|����t�.�פ�0fMJ��\���&$ǔ�ͱ��}������#���jA�H��<���㇗������6�x�,�dp�ވU���1���~_H�"�5Ѝ�*:�a�������=øޛ�Y�b�<���iF_���JsO<Q����WӋ��K�/���Θ�GI�i��3�5�L�<�W�D��3��	��l[Җ1M'���Y�5�l`�^����J��,o�1�`��̘���e(�D�TE0A��[��l��SVS�x&�C@��f|�u��.��<R��/����R��~�F=Wާ��+oȲIG�8���qᗏC2��Gϯ��~�'ב/:���Bgw'�&A�k�E��P+d�W�N�БN	�&�C
�T�E0�������hJ����(��� e��T: gL�e|�����G��t�)%z������\���ewwO�� ��9W�$L�Znk���e$�k{y8�����Y������Q���6�#)��q���ٷ���@m�} �v�Q�M�	�w�k�"72(Y��'�����Щ	Ϣ@�LMG ����o�Q�O/C�D�\ÜY�q�׾�]gs�Q��Qw�����X/L�d�:�HyȤX7.#xBh�Fћn�'?�{��k�%����)�1a�X����� �5(� ���h\$�ܨ:�it�Ӽ�X�&��o�}�U2`�|�||��c�VB�&D�q�_^�s�W	c��e���HG��,�-¾:�"~p�Y8l�d��Ƀ�X,b��M�:e
�4f13Z��C�<�r�{Ά̓x�EX��f�|�#l�>����^�-\p�q�2������0_>����L�:R�H�#�ۨ �Dnt��}��Ͼ�)�j�č����uk$�a�]wӹ�)�K�����G��5��g�eoa��0�9�G	F:��������2L��X^9����W�����h<�P���� ��kkFΔ�����7-;������$;q*�"<��zsS�{%�r2c�"��@4�D��z)��0���V�W��fƔ.q6.��4b\Lw�d�6b��2���d���s��4s%4KU�vzI,�YvI։��Ӑ��х�Ҥ�3�������+�-�~<����=��kw>�GMf��H%�8���k���	c�`���U#��z#e:�DD�e~͏jEŕ��-?�W�:���*/����5�غ+^{t ƌ��f�J�r�jES4O"    IDAT�_>��(P�`�Gc<`���{o5����\�f�熲��7;2a�Q�(��RU$�+?�/,C��b�������OS�[Fɘ�Ӻ�ɮn���R�.Ӎ��01;��mqj��J״+n�Ԭ���4Fܓ��!"����87�Ϸc
�ih���?�gɵ��.q`��%ş]q�H7�ܝ�����ra1��X+�3�ۼ7m*؍�U4�8�S)�y��l�4ͳO��[2K�4��<�@m��.8��Kyv\�)�,�d�2��\x��
~��ǰt�F�C�@��ݠ	P���7�����H-�J%J����P�s����m�k�����ޙ�B��mӝ�k3��,.	v�z�6.贩kS$�?���Үs4Bʭ+�*�L�*���Uh�Fa�+�6� �h8�x4"���T�4�����(�d5��M�1�$���JM$��r�RE3�XB��J��'6Ȥ:�J�Ŋ?"��&�z_H@)� $�3�	���b��ys�m Gv)�PU�H@i�>��]2My�,h��m��m7��V���ұ��h	tFY'�tIQn(k�.����P��'�r��؃n���F&x����(W�<�*_�Cy�N���3�802�<�ioj9��sE�_�15����U�nO}ېjE��3��Y������S�U��~���sy>����?x�-|�[�a0��5�f�%�Z��&a��QIF�v��R`:-!*� k���Ǹ�׋q�����E�B�V|U�}y��k��w�����s��	L?�
\����O���"�r�n36�g[HTCN 4@˿P��}���E��<�Ƥ��`����5��v+e-��@�S-d��c~�S���L0������
.��0Bu�=�Q�Ѡ��d�XR��Ui2��u(%e��@n�0
�q�%���
0c*�2FR���qq@���@=�Cn� je�q2�4?�Ѥf(�>�;�L��2�b����5M=��p�A3q�%�I�69��6�e����>���ߒܽ�x��/.<�x$
L�Y�?��Ȍ6�/��ӇdG
�	��k4��I����Q-í��'����͂AfU�fa�`� x���I���V����I]��yg�K�;:�(�����?�5��C2���  n`Lg�~�Hy;�a$�aV�����������NG�۬	"��/J8��h��;���7� $�e\=��<��j� )�H���i?&�%љ#�!䖅I>��C1e�D�fo	z���7�&y�UK_� ��x�ױes>�m�*����M���K��\�݁���0:���&%����D��"Hj��E4P��_�'5c{���mêw���K���M&�Hw$�ps�9 ߏ���0X�~#��s.�8�d���b�~~�X��FY0G����N[�
|�n�=�~�u��<��&W����\�*�!���2�+/9'5	����\.W�Ƹ�cD����%��bN�)[Z��׿y��5���?�Ǟx�F�_z����j��cX*�X�'�7Ѕl��t��Haɩ��� �����.��{c������s3��\*`�ĉ"�j�B+�l����a$[Ŋ�>���a�hU��U��x,�/̛������YEc�*���������[�0�mE&�g@��M���u�N�l�
�-0�i��)�Sn���� �6�Cn(#Ns�T
�1}���hn�N��A�k�ds�ET�FQ����*��]i��Rpc~�إ5O2��F�Q1�pպ S2��0E*=UK�!n咲����3������3�1�������+;���o�?>��۲�T�p��� �C�톫�u1�M+��t�����@�����D�T*T�9�ɟ������h�:�c9^����	0=昣��۩r�]�����DQq�����+X�TڮE&e���z��a���B �]а�Ɖ��U��7���'��1��[q����,�xa�8���y̾��0�#�w��/��N���' ��װ���μ6��ځ���`�2"���#�l� ������|"+m�ހ�wj�eϭ�"(���YM��X�,��PLZ�K�fJ#K�v�e�G�b�I���z����[�s�*)�Tp�r��"US��Cl��� ���߁[����F�z�|ܡ�:.�0�
���릡�v ��#K��ka`ąHʘ�[e��,YEc�bUCܹ����ݪ0J�b�-��s�6,���	�o�>V
l�Ew��T���p��H���X�))��,���f��5���V�ʫ�^g��"F1�5jI�7��DO
p��VXm [�bct��$�]���\Bv���_k�tS�X7:�k3]1�� �f�2>,(E� ����|�a�l _��aeI�`0��fk����ƘK��EvW6��37,Ϲy�	|	�XS�N�\�F��&�O4��M�0Ϻ��2p�Yt��}�����c����R)*�7��q��.���V���QkF�������Ha�xb���񰐎K��b�\�#�j(�����g0d�J�����F�^!����{{�Y��M��`�f���}��A2�h �Ǌ{%j��Q3L���Mf���P/a׉)�������z��y�n��U����PE
U*��*@��YS;��+��ч솴ɽ����A�������D?BѤ S��1���&sY�tG	���I����V�s�{'�jy�uY�e����B���,���LR�I��˹�J�iX]y#A�D�T�5�2�.�Q��8TG��2�T�$6G(�9�5*�̌hK�5@g2!1o������.�da�J�c�օdte����Y�� ����j�mC2cJP-R�hX�i�aL-2R^�9�ܱ�1�+�2cZ/	0�+�I_���.>�0����_�(2��q,^�.j��!�v����Y�!F`
੥������h�r}c�O%��FM�,Z�������-R\)pDM[(���QO����%�{1$1X�q���i�p_;�\r��HG�m����ưHyKUnaY|���4��F:�>�g'oJC�o(#�l݀��)��Wb��9l�R�f����KV~.l,�p#Ѱ	���]��Q+ �RSM�xNy�`����T|����I�9�"6�_�7$-K��@5��v`/-�]��j#�Q(�Qe�S��nV"W��&�9�c�]N=6� �_����%�!��*#�cҘ$&�q˦رm+��[8�2����C"�[�� �إ��F�%�2mN:����/���z/>Y?�"��C.f�2	����Dc�5[����rm	�%5J�F� �
S�)�f2�<��@-�ys'��ӎ��q���Α�p+%�2m��7I%Z̆�!�����@�PG��_7��v9珘 ~�����4�P&�k������O����X� �#� &��A���!����>G����F712��H���;q
�|�fi��qݦ�x���Pt"x��WP����Ĝ����+��~�;֮��[����`M�t"k�Rk����ΐH�,��Z������iK��䘦�O�Ѡ�Uf*���m2�>���1-�d��Ǹ�x?��a8���k��:�%�W�2�Z`���L!L�(�[n{vƔ�)��2*)[ÜV�cD�/�i��A�%]�6ؠi�}�;$���:��I�1ّ��ŗ���W���Ј��X"�)������~swE<�Ng�	<��g����L#���0�jբ �c��߾�]'*c*.�mL�l��ٰvV�\���>
�=i)uB����c`�zD#��D��<��\��f��*Z�m܂�q����0U�H��F�^\���+N=�t{�qҔTfKg�_�(�ǟ_�R������c�Ø����FȘގ�_� R^S:*R6�5'μ�TȽM��wx�,�+��(�V�eA�t����d��4�Ζ�L�)���Ah���d�'��@�jL������z�<�/�sj�xy��7�1��d�y�7\%מ<�����wR�Ł�oh����i�&�{�������[�:x;i�+D�Y|q��Ҹ��k�4��6I+��L�2��xv>��*�����2҄/����S�����ɜ�5\1���Hޗ� ��Jć�5j��V��8OP��n^c��"�����V�óF5{�,aP5oVOT�/u��&�0�}�/U��"��H�'smZ��U�AU��-���1143@�{�z/-h׷��M�$��6`�ܬYU�,�����M/{���i|�]?ڀ�g���������hi�Ş���+��۞qm�z�gM������$ٕV�#�W�H�d�+�
��Q�:�)c#8��q��aL��	�
�A�JE	J�6������W ���X[��"��sC�� |�i���ܠu%ng�=�20mB�w�T��}��ʶ��a����`YV������|�����f��ʎ19��q��9m+%�n�->�{�����8�]'$���_�=�%���U�����a<��rl�J$Q�ZA�^F8���&����n�z<@^6�82p�#/��o���,!	�X*J�GM��ث\m�J��J N ��1��P`*o~��4�ox����FU�VQ�Z�W�F��!/$Δ�~�����8�%Ղ��(�b~?R���ʙQ�1)/�t�MwJdK�/�Jf�C�?��n*S]�C(fr�V����Tʫ�/>��ѲNׂ�ń�*0͢��+6��aD�~�E%.������yG�Q�z����-92E��������S��R^Θn+4����{B�vF8���p�'�, %ZO.���܃�Q�*�?v,b�hH��t̸pe��~T�cSC��gg��(�B�t��/�1����
) ������|}ϭ؎���6��	�Cbv�a�m.�JN�$]=R��(�B�BM��d��k��|��y�F�tn{`	^^��d�R���ue(����ZT��5j��Q�mE�Aw�������y$��;�[Ui���xh���)H���rU���Z��sl����Q*��L��M׸�!k_J-���3��=�n+�ޟ���n�a;�,���s�e��*J�2'v̑bϹ����*��A��"Wu�epۇ�H�z������{,V�	�,X���
�� 9�u�Qf��&|�-��� ɮO@cx��!�1���BI�v54k�LׁD�Ew�P��(N<�P~ȁ-#)bgL�F���@浒.Am��ђ<����^�BA��t���|	sf��x��,^{�S|��V����`w*�yt�8�z��Z%T38��p�����'�`��=UlZ�sfOCW�Ѥ�L��*[�DH`��r�e�}��S^��C���q�E_�^s�dV�A��.Z�{Y��bP\�≄��:C��
R���a;ar�$CZ�P�C�}-`�]!��g]dx���ѐ��1-�:���n Ny�9&��x���*��4�4�a~1?���7L>G:�M��̘��/�;hd)�-��W?]sL�l�=���9�i��L�#>2�n��6�������@���C/[C._�����N�Й�˽�kb�Ni��{�=��Hj�ϏH8�B>�J5����i�>�"F��[�h1ȅ�n�:Q6~�����=��>Ji�����RDBA�l�	��%M��yb���Ø8u��{���)L���^��˸��{1m�\}��H�Tr���Iܷ>)��Ͻ�r��YS��̣���N6��h���ߎE���L~�ڙ{�Oh�|����/M#ð�-)��Ӱ2Z�����M�������x �)U��*�u]��(���
(�۩4�����`��4o��[�����J�n��=����ޥx��7v�M�7o־����ʬ�\��z�"W�=��<��m�9y�6�ߺ�v��%�1���0n����2�bU���0>X;,���H�p\�b��v���mr�̲�:�T��ۖT-	� f��M��;�k��gFcw<E����ֆ��&��8����ki6�Vl�Ja_Kk��'*}��{��1�)�͍�
�֍��k�Wɺ�给=��)����B@�䍾��,����
�mS�A���Ǩ�2�X�ރ}
�٫��ak��h3Ļ��$4;�'�o�,�jZ���ct� P&ZH�f�b��ճ�g�q��'a�SEU$��z��W���^k��q�c��«c�D#���V�E��a���|=�?�z�o����i����P@#M8i�+ U�^�g�L���^�:��u��oAR��-_cb��dY�\�}B�-e���Fk�ɨ}�5y�0�ڬ�Bk��b��7ʨ���%�t��1s�=]��73�f����ذ�4�S� �Ҕ�꽒gO��&f0���*�&�v U�K-gT�qL/_���Ģw���p�	8M�!�t�H����TE
0�=�k`J穕��r&n;G,0��E6�q-��Q�9
��5��Z��4
!B!�hլ���F����Hq�g@�w�ɍ�B��H#�X`��)�(�%cJƵ.2j��=�9����L�H���0�dL#�����Y5_M���j �=G���!(`�3������?S2��r����t���:_\t����+[�������3V$�N�F	d����|�L��`�]��M�Z�N�о�ْ�,���x	$k@=��p�y$.:�0��ޖ��W6�{?�ut��Ņ֏'������pЩ�Jo8�©2>�(����p���{W����ގ�;�{	+W��/�D��p,L;�jv��
��O2z9��A��h��࠽��kg����EB�)��Ư���hFd�\�c�p=��W|
�?�r~_JdД���眈Jô�~�B:�����^�6 �HH�[�Z"D�׋����y��2
C1�?��=�B�l�E'χ��"W�c��!��4�R�/׭PjH��9T*{���}C���h:S2����F�fK����D��YY��A��"��¾*�vEpͷ/�ч�,�Iȟ��F��Z�3�X��z��똀�_��^Z��e�=]H��r������ñ��n��<�H�d���Ҩ��K\��I �)\F$�bڤ^\q�y��!ı���O�D��n�����;4ZÖ�
�~<��R�|g5�2�H��8`�ݰ��itL���mA4�#�^[[`���������++�Q�����U|M��1U)/��t�8YAc!mGM5G̋�1u�Fz��OD���G�ɘ��"G��2��1)���!0�tI�i=ܔS~=�)-ֹw�ϗ�X~�ZȌ)��\�|n����)�J����1�Ω�H�>
�Z�1��w"fO�"A�ݶJ�눏�A�,'�[�����;�~
�ˡHHt�)
\��"�<f����]�Y���*+њ���O��׬���C���Kc�A��Ê�K�BKy~�8�(�&Pc���d�}A�`̄��c�y���U0v�\�K�,�m�߉X"��~=�O�3	�O|x���Ӛ��S���b\��
��׸�kn�b���0��>8ָĜ�R��
)�dQA߄e���A�z��b
�����H �El�Y��8��B+X��b�t����jZ3Y���-�S��֜��68K�LB�����ԯ1���um��v�bX�6f�~T�xMf�쫭96�$jQ��^M�|�L7����؜i���sp�4K;06�ĕ�<���Gs�)u��y&��,�̚������C�(�H I�/�^ca-�%��f�꽶�o���S�[#)�y��-W_(UʫϺw_-;.�T��є�lE���מ�k>n�-�B�b�'9����̧>��I�-�4�<�QӾoe6��f>��` ����:�zZh��^_�l�����M�Z/�`��j�i�O��g£ωIr�Y)d[4���0�s�X ���U�>&L�I��\2$�L�{	n9��t��C���+.�2�����Y{��'��b�S4�O6TpǽO�w�#�Dᆒ��b�I���F�    IDAT��T_�T�
�tד�{׻��2W�:�*���k�������l�M�����"_�p�j��5+ܲ��;�6��Ei��DڹvSx� S���26��YԦ?k]F��n	�F{������v�����C@j'~������[�A�6�e5l�J��}�۷\2W,[�b`� �Q�/o{�j�O6�`�MWGx�+�4�1�k-}iH�U�Y,��@�0�\�l�D"�`�&�4cJ?�6�c?������%��FC
L;��������ȩ�1%0�{�4'#��!�A�b�d�zMß��Qu$��Q�59f�N�k�3����ښ�¢*(% %0�l���G�,N>x�Hyeƴ�6��㿏4���9���1,}�=9��A�&3�'��ӭ����H��R͇����%��"0� =܍~��r�L���°Z�/ݼTj�����k%��]�b�e�����E�Η�0��{��M����@�I�Fc�h�DJ@�C�JS��b��t���`���[�|̙����S�Ą�=(�ز-��KVah��P4-U|�R�4xp���W����P�~�=�8F���7�_9�`��t��y�M�M��yP��E�y���yO/zu��?ԏp�>Ju����k��`�?�`U��u�4EehV�iD�e��e,���WF.(qVs��n�Į .9���sv�&���G�m�Ҁ Ѝ|��V�������}"I�T�&���*F���ub�a���l�`;U*m�O�u#��)m��ք�9ED��wp�����"Iwn�bM��f���6\ï~����&��435Ԙ�e֤J-[L
e�� !���kPg�8���J�[�4٤(�P-�P(���70o�t���1�/֦0�Ҹ�+y6x�(#�d���)���s˰n�b���ģ~t�����Id����H]��)N�nXr`i��ExE�U�G��@�t�O��ӌ�Q`J���,�����_���mЫu��ʘ��1���dX�42���#h�i�PƔ����E��K�bja������L���ߓ�	�+�W���mS���^��x3o�la�)��Y�SEe��L�~�!�uZ:8ӫثU���Ǫ�
�*��M<��
,Y�!��4Qa�h&�_4Q�iė��1~���0k|�+R �Ǯ��L��lX��z������i����g�|�B.+�C^�h8"�}�H�K�aʪu��,��O��sۀ�9@��^^���q��~uӯ0qb�)Y��_����>��̘���c�����(���aђ���M��To���*�0l�e�L�걆ҵ��O�15�Z��0�^�m�<aL��`��a�,��k"�\䠭��\y���>C�?�%E��De@ĵVd�Q�6k\a�4,6�n��m�B�'��R�ɶ@5���(���U��l
�0UYa��9L �3�F�%̟*�B�&*����� &��p��G��WpjfN5�˨�h$C��A����CO����Fz�c6x �`$*�^�W��i�M�����\MX)�� �%�3�ـ@���-u׳F���!'���+d����
1Y���i�sWy��s�3��W��6����ܬaao�-��kf��Z��o[T��W���1��ׂ�{��^J}�,�M�����x���lE��fO��U��{R������)0,�nd�f����ys��+;�璲Rs5�~U���(�l^n9_-����t�!8���0sJDw��h��r(eF���zPF+�ۊ��`��4���\!���ʔm��4w۲�m÷�0W�4����&�a����}�oc�[wی���mҊ �����O��*��T�X[@mׇ9'쨃���o���+�ianeHrܯ��|L����`��ˮU�Y�^�u��5��/UU��p\�E]���¬G�82�T��~,xs?��^���h�#-�f4Β�ϙc�OT�&���x
{>�����fy����,aL#a�(��/��N�2��w�@�4
0�dr��h�UE_���4��Έ�/��$����Z=?�rC�S��d�	'b~�Q�KE�S��;����G*�29�1�y���h��E��U�l�6����Q�W.hI� *|���`:W]|��n˹��]0��L�8r�~����/o�Oo�2*��c�!OHL�)�q���0eow�[�R����)��n�U6���ij���3�̮��cq�Y� �9
L}i~|��Qr	L#��0~��d�i:Cv��?fa3VAXO�
�	�yAK�\tv$�EPw\�����PP9�Y����l-hR*Hj�?�enb��6D�0o�^�s
g�vAӭ�}�FN)�4,ΛaE�
>���%���ː�t!���P��@Lq�%W}��;�9-��h$�����X�	�2�T�̽�D'.�&|���r�o c;���;_��=$����+P��ϣ�40Zt0��,���	;r�(�z�_Q�:����_�	�"��F�$���N��O:���T��n�+��GjV�
;HGj�p���z����nv�k�g���`�����U�@���/�?G4��r����p���f]j1����d~iz�.�H_VKE���a-�)���3�pǯ��cb��񦽼����zSWN���s����`밋m��Ov�Yc}�����e�����G�/��}�k��>vjw�ŒF���2���������S�1�D���	�u<W>W�!�gS�W�U�;�H��`Z2.ƬY��P	�6����48�j�$�e1L�0͏�٥d/Q���JP*�.��\I ��Hy��X`Jp�~Z�ʂYs|�N�
�F�60ml7fL�þ{�������z�{0GE��`0���H�f���@gW��q�q&,�b1�j5�
�p��9>"Fl:������{���l�{ﾏ��Ag7��6���[�	6oBgGZ\�9Oj�7bqu��ۺm;����I�0s�����ߔ	<�ju,x�%�{��D��7`��-�ͬ��b�=��*������'9��PB�wE�Ƞb�QGFgt���OǱ��:����tB%� ����~�����{������f�ˁ$'o���ϳ��fKw=�LX%��M�G�9�uwt��Ư�
˟]�Z�g�B�g�8�
�ޯ�L���mf�$�언� ���Nw���d����윲G@���I���8`����T�ͨ2��mp�����G�Є�;q�����=:�ԨZ�T�6$�3�s(����C���,�U�|��8���*�]9��#�-��La��6y.W�ȍ�B�2��v��O��;�)���f�+松�n7�� �lA'����f4=��{��"���[��[fT�
o7Qr�_7y�9��"RpiN��pٹ�qE/N�ğj���R�� ����5H*��9��.S^˚�:��W�~[` j=���Ń@��s��Ѧ+2���@�M����9Ц��b���jYfdvE��������ۣD�jTm�[�^_[�&�ڐQ:��{Lfg�3�����yI݈:J�1�
CWG�p�D\���q�	�aJOH��pvϢ�ۙ>�����X���J�d@1�2��<d hQ���}huӖg���r��ޭ5�^ޓ`�г[�S��6�j���։釾�kb���/���TМv���UO��~,�9YGJ슲�db֬���QW�o~�#�?S�2��w�~���9iFj���d-m�]�;ۧ�F
=ܭ_�3���6ex5�����;�[���׉f����x����:��i��)�R��K��ݠG��i�P(C�-%�4И6����7C��4<&�G4���UO6Ib�����0e]̉)�iԀi�:U����;�шEQ�(0�u�W�8(��-G&��s�+54��::tb���ZN��r��>���5����Zj�i��C{h\rL�r��".f��=�5���)�4�ʴ �sEtL��=Omſ��w+�E��7e�hL95cg9F�a�� u���bHE��8�A:|r������gͻ�)�iu�2n��|�#'	0�b 0�g�f��&��iDX�g��"��ŋF���9�	������g��1D*oM S"�p�Nt�}g�5��R[�(��0z׋�zD*{��m��:q�%�cɡ�|J)�_;~$Y {�X�0T��?��|��ĒSOt"N!�	�Ӧ4���ѽ�Z����;�R���Z ɵgF�m.�
m��QفI�!|�c����*���:{E¨5(T*h�Sؾ��'W�����)��z=�D�Ml��Rl�M������B�u�jw�N{��шI�:��p��- ܨ"�,!��#Yŗ��*�p�|�8+�ĵ���-�Hm�HN�W��k<��z��)�R�� :^�쫌! ��h���tZ'�QH`*�iJ�fl�tt	��Qa|Gi��>,:����?b���ۺ�J��9.�>���#�ͷ=��߷�Ƙ�0�x;"��9)Z�������FAwT1�
�Z�-�����K`�OL�P��hL�=hK���2P�>�{�%͏B����)�R,!�ގ�)��LB\�Q��W�F�kѧ���J7S+���K`tw��&"Bo�fͦ��gb�o��Sm���G�2�5`�
C��՜�ɎF
E�*�<P+�42�fq�F���L��H5��`�`�\A��@�9��$�X"m�H�u"*M�$�4U"�9Dì1����Λ����oq@_̺̮ ��J�q׮=X��:y�bt��HK���7+�-&f{0��S�M�|Sˇ�D�v�a۶����Lìy՘Ig�o��U<�l~�[���ķ��-L�޷0}{kw?��r��K�:ڕzWC� 7~��X���B�8c6��e����i��y�E�7\���i�$����IP���!G��\��~�M}����i�4:l=�7U?-��S�S�T�`*%�v��2�/�Z��X	k�M�Z��{}��ttS�쀦/����G�V ��Oc3)`��V�T%Z��He�a���}8��hV���#���W�����lL�$ʦS���^�ȠF�&`�v���Y,{����&�$�.�=rd�$P��<�tD%Cr���ЧX�Z>+}}�0��~�y�R�j9�d`j4��ɵ��i��4��r�ڽ�5�/��Z{#t� D轓5kF@�4�:���	��li��	�	ֽ��W���Bͦ<r���r.��<O��iQ�5u��M^%����A�w�{��,^�*PuIʜ�g�4>k@�6r�r�Y-���Z	��8�QL�N��c�S�D"�Q�_�f�:E~j�ǁǟ[�_�M��Ri�Ѥ���ͩ�6�=��#Hh�� SӚ7�}��&�<����zK|���{eO��Ѻ��C��wK��5>]�/70�ߖ�O�]#��a��Z|��A��2y�c�!~�HC���*n��L�w�BaT�A h��`v������S���@�]J�������k����K�p�����0��iTQa�	_��k�&'��4���[��Ŭ0U�'����71H4�x{F4�^4�*�J���/�z���mQu��ĔT^~���S���+4v���Ed�L8,�4�A&�9��r�%���2��1��'ߺ^G2�k:FihT�)������Չ��N3*o�r7�7T�(]]*ɋk�i�2��PGW�K01�?�:`��[���^C&�Eo[��v���A롻�؄���+FE�8e�4�S)5<��T�s��Tu	�����\T9k ��-��Dó0�bCn49�e�>�l\��'�8	�M����'7⟿�tO#pK����B��Y�r㔎9Y8��8+�`�']�N\��s���t�_)va�(��m���0-�A{c;�ŕ���8���̩��uj�ĉ2�x4��|xx���*�K!���d�G��%"o�����u��b�֮�u����7͜A���E@#��.�#�~���>u�e8��CQa�<_D�TA2��)/�~��;�qߟ��+onA<�q�jԤ�vkXt���uX��ko��qT �Ms_m�I?�ë���#�@&Zė?�Q�r�BqW+s�3�N�l�v�3@��Z_��mx�7Pi�!�ރ��^�J3ˍ�)��m�΋�T�@�cQ�b��ij�eZϟ��P+�Z��8hV;������3�]r�n-Z�Y�Ȳ�&�/o���\�Y4�YĒ�Ҁ!�qńt��4]ׇ��i��]
u�z=tB�T]�21���6멑P�#����p�X;�-(,� \��6<�����*2�6�ʊ!�j��C��8ʣ� H���F�(U>KA�J!�ݎXgu�'q�V�w�>�����10E�k�^ՑR�9�c��?d���ɻP��_�H�X�ax�q�G�`�:bQϣ���DT�LG7���HwM�� eS�C���&��hR�����"����
f�2ʚ^��	
X}�J�"v�ރ��>d�,C�&����F�!q1N��Dݨ�ґG�}��ݳ��NǴY�)�N-��"(*X��9������ \�+��X$�R�����^.ӅN�%grbJ G�@[G�/�WX��:�C��4k.ڨ1P�n��WM�먧�,Q�k��%;0 ����(Q�����6���}�g�3��Km�R�u�	4W�W�ΡW/����Rkp�(}M�gZhŊ��x�1�-e0����sD�(b���eZh�n� ͧ����~��=ѝiN6AP(�&��JCYG���F�����rH{�s��z�i8dn���j�2�I��#y`ŋ[q����M�h�{Q�(bɔ4��\j�� �%�b�i�L�ײv��"�S���(��`҆��B���$��d/�{��%8+�{��3�1�lն�2��&�Z��>m�-6��lrZVݣ������� B�:�s�mc�)~���ʃ�`�.����D�o��9L0m����y�ǻ56�3��h�nz��d}2���k��)�}&�P��j�%�2�jU�*0	���*�:t:.>�X�|�A�nW�災��Xu�gT�����S/���נ�D�K����R�:���!��7�uɞaͻ���}�3F������iiR���4�[��O9
��TL��w6�w篱�UYW����Gv�����V�ZsK֗V��g��&�����,S5Bj�^�
��VC"Tƌ��u�b�p�����%�����J*�g�����f�oDA�����D :#�+"�#a����w�竍��:��eO?�6��`�e��(��1֦AC����������C�̺��VN
�N	iS1�����Ry���9lFN�S�������4W@�KL;:�LF�O��rd�ɐLo>Ѩ$B�f��H��\W�v�*���S�Gl�k4��ޑL"�db[0�#Ґm4?J
����������T��t�T����؞�7P��8��8.`����`�w���r���:��6�KO?�_�T^ w=�	����+�P�E0m���E¨��"P&J'U��4i��Xn4!$�{�@�a+ƥǩ������5�U���Й��=���D1�VFw>���﷠TO�&���{&H��l�W�n��:n��Uf����)���	L���P�e�ת�zp�h�D
v�]�K�}��H3�pi�C{p�������`�t��V�@ ��&sB��x�����0X�"���H���Uu�t���e9$�#货��M�:Or8�.�)�M�t�G�)1�YA�8���6L�
���G.>�#���F�ZC���1�RI��M�@����}+_~�D��#�H�=�)� �Ah/f4�4bG������e�Mz���Jc��Z����ūp�Gplg�ԍ���T%�v�8�!0�ֿߋ{��*��,2m��vvE���	���i�y�h�/�-z4I��5��f5:�.�v�<j�~<�?�����E6z�^�����2��<��������6H[�����s��Pm2�L�͋�]��T�sI~^W_p���Z�<?=r����,�)�\�N9�L����Mc:8�z�*�G]�L��D�o��a)��$�=�	n�    IDAT��������ށ���,jQO��${Ψ��;�YD���hK1^�#��4>L]A�k��s4S�ↅPY�_�X�ʣh��,��,��O�76�R�4ڲ��v��{�̙w &M��F,�7�}�5�wa��@4���g.��h��5Fq��~��/cz7D��ni���҂��/��-N�|��|IS�^��Ш�a�T�4�:t��r��޻w�lټ3f�´Ys5_Z�Z�%#��Y��=ݘ>�q۵u�S'���"���r��4�q8����ŕw�9���S��C����9 ��+g��LY����M���1�#���t�Ll�,b��M��}��;�u�'��-�?��j��|إn�\���e�FK��֖{�[���11�XkCN��P��t��&;���J�ӊz����C7]S��z�u\�x~^~Wgj��M�b�i�g����8B�!,�Ӄ+�?�z(:���m�C���G�Ldx+���7���e�8��4�EĹ:�I���cFt����vL�=a��{�})����=Y7�����͵�n����&[�������\� M>���2ja�'� ��g2��k:&��+I�3껺Ƌ�V+��7m�Xq/�o�/�;�22!^٭� @$�s���]wyjj�j��Z�j��������A)'��N���h6�e�R#;�ZA�0��z��gM�G.:g��3&��������#ZRN�7m/��o`��7�i�F�Q�ҽ���5����J��g�����_[�@hskI�E�m�+���V˂�B�)�i�[�f��Rנpu���ӊ����ێ�3<�94�����?
� 4@˿���֛.9��6�$�I]��=x��^QR�Fљ�1e2TE�.ߍ�ԟ�r�g�	ࢃ�}���5��u�ф6(icC�2�Z�촺�b��<W��W�a4�	�X����g��e��Y����(��t����s���\rUW�"�0Muv"��;����,��H�H`0��tbZ��V�%�G�L�P7�r(i�5N*��8:ذo�Ɣ	��`�%ìK��".6�Nte�H:I���)��rPok�&��*�K&c谹�LT����'�謚�B�q�5�p����?������h �ď{��\�x4��L���Dr�hω�]�m¿�t;�+q�HM�1C4�21]����w���14_@�o�M�fL��2�d^e*%y��9�mU�pI7�s��ՙcZ§�=��D�I&��B��������f���f�޸��K�^�p�n�f@�2WB��L$4�Qt
�/Ʈ�MT�c躇����7��9}��>�PI{;�PC����!�ctb*�>Ф=����o\$1T�p�c����=�)�3�杈'�Eߨ9Z�:����̺�A��]�B������Jj�����`��[��Fi��]��ŗ�x=�,��bq۶�Ħ��P,��i�`b�DL�=�p|��Z��9n �c�ip�R*�zG�g'ؓ���
�7��Gic��C��ټ�����0��+��?��u8�ňH�N\�C7~�^q��0^%0�>�&r�8�;{��;I̤$�Bǩ����e�+�Y#|�kH����R3	�b7�����x�$|��|��8��GɃA��N�)���o�n��TЅJ3�T{�8#�3)5��)��T2���z۵�w�5g-�M�\7V��	u��0bm�:�ҳ�?�H��ha�J�nA�i��>��R3!SY�6��A�."���U��V�t���6�S:ű�� A��ҭ��0��r͏J�Vӵ&.�l2��#�����Q!V>#�J��p��Kp؁}�J�#�XDk$�.���<,�8ҙ4:�����;p�]+0\!�L��H(05T�cL�OM�g��;L��=W��C����',���y̴�Ia��K��Ğ]{����w�D��N@<�@,��a�s��]شq=fϙ��(9��Y���a���h�tQHh� 5�����y���gA�<睲 =Ԙ�t�
0���өsB��ul��-tnݠ�tN�:�֛�i�2��ٞg����݌�l�S�`"�&��Z�QI�$����xJ��Q��3�kL]��!�V (`�&0�Z3ed��ML��=m��dY�֞�H����^�nV��v�T�ry[����4E�
q��i0p�3+k��6EU�EH��Fn��8�=a!�xÕ�35�4`k��Ϛ}q�,�l����W��G_�h��Z�)��n�@�=+9��+H�cf�LS\�#{��͞K�_n����^�DO�1ރ��ZW�q娰�U�cT�,���-c���\�!$n�Q�ɡ�d�L�ݺc�0�5\��=B�w�'��3��?�����k�@���\��R�?e��:ҿ����C�Z��������":鷽J��jf�Đ@��6u��*t�.�#TEg��sO[�+.>�<A���������(W�m�/n�/���Z�T���8�r?�{Υx絕���(���H�x!e1�6��^�a������tsϞL���Ё�^�=i�3�S�~M��^?���kFZ3&����[֬�����q��Q���ݹO��zV�ԑ���Hdc��1�
��hT�Q����AW�D*q݉S,�&�j2V�M���/��hғ�K�������>���/�=�I�"�w n4��q�rj�Hv��e��#g��2(�-��84�}&�.�`��]SN��
N���l"
	0��Ɣ�x�rM�7�)�U��0��:$^�V����Iʯ����0��4{�� 4?�,�8*!2��+DTi>0��� ��`�T*/5���	%-�4�T^Y�<��� ��w�,�j�z��.9�`�ç�9���,?��}x�ٗ�$ћ�㊳���9W͏<Ry7�{?�#�
U`����j�R*«VQ�Q���|^�*�T�YTD��R;c���	A(�)$S4�Qp�~��i�e�1����-Z�箻 �]v�LLycK�Om�?����lG	D34?�h�n��b��F�*�C�D�I�&�He�,cqJEqv������H�n| L�#���W#=X).�0)U���	�
�*ÈT����Yi\|�X�h��F��F�m���d���\�7�«��Ŷ}a���� Dc����h�L���_�O1C��j7��b��#�b2S>������Ì�ɣYCqx;fN��k_�4N;�h$a��5�޵;v�@�HƑj�F)��+^�ko����"<N�c��VJ�l�F��rG�-�t�k��/�� �������#Zf���4.���+��?}��}�b�!g��@�#��U/��2���?�[�x�z]��;I���ŷX($�$�q*�% ��,�C9�����a�)�#\�q�������������D�@<�
LI�����{����U3b����Y�5�SSӥXm��wl�0�H�?�8
��Z��"��511?���ִk~��˾@��@}4�u�*���N�$4�J�)�TrcH�(%�<��(��Z(��	0MtS�OCNL-�֒dBr�&-�T\\�П4.��'���L�3U�K1QGo���˧q�t�)�����u^��F��Og�Z(���V��o~��4��tfS�\E�6��S��o�4��(�CZ ��#�$��ѳ����/�WWˇ:���0c�tL�҇�ּ���~�dUǓ��2u
2�4ڳY1w��F1yr�Xr$&N�$����q����î�;p��W‹�(�����RxsC�<�$��p�����#�W�v�L�'���z�S��`*p�i��[���/y���b��MX|�M��߷.�S)���ud�� ��_���]�
��O��KwX�j�`?

����~�Ci��w�/�Ѵ�n@�X#,Pyn)F���:�ґ�$���o��׊I)��^�s�.[�����N�X�m.:��)��K�lzf�����Kz!��x?j��p��}��5��ӎBWV�+�YfSL��H�
�
�ࣛ�~�m{tz�KR��HvtHF9�D</�]��>�7���d��;wZi�FG5����H*������������$
��� J��#���R��$OK�ؤ��+��?\�	��_�R���j�����@�:��/� ��_yi=��s�����˝w�ױ7����[#�c�	|k	3z��Nr�:��b[�6���(�r��۬�Q+!��ȅ3��7\�%�z$:�i�r����B�
��������w<�����u �b�n^T�`ԋ�����,�U��1�3G�5�&T�����M���]km8�}�3ϯ�9]�^��`��ӺcH��3��L\���s�z�����h�����:���������g�]�]R�f|�Y��>+��b��L*��Q�����F�ݞDogmmH�Yʤs?���r�J���\C����R��&{0̨A������Ж
�=EWGJ^�\����B�E�Jf����=��O���zm�
���3�Ѩ�+�f�<�	L��H� ӄLI1*��<6eb�%l��1�s%��Я7�Ļ:D#Z��ēszY��h ���?��RK�Ͱf��/�fB�NQ�ȺԜ�e��ߏF��cL�-�T����M
��֜t]7�c�g"ٱ���KKD�$T�Z��.=��=͏�j�H/Z֮�kӑ2��[��c+^B8�@o6���s,��s���G*�f|�wa(B����S���׫���
�s�-�4��&Ø2�S&N@[:#��|Q��}� Fs4Ť(+�4��%�����3�ư0[����jV�^s��>0��ѝ��Ƿ~p+���df� �fP,�P��Q+��Ʌ_�����+ 9��J���� J���Jsч���r%9��I��HqjV�b)�>^��d�z�� f��p�����A�a�A+h������T*(֚ظ�Ͼ�>J����`��q����	���NCni��-32���AR�H7"N�ٍ�JoT��LJ"�R�q���T��4�o|�s8�����o)|j�:*�*�^�G+���X��F��/����*��-�I�=�jE����l^Gf��*��$�I���!��D�$�X8�R~��8�<�%|�?��OX`y��Va���?��1�U����#���0^�!�>�O�U?i�$�Ձ54nHl��{�W�{:��,z��¡:�l��q���_�:3<�5����MK���g��<������`��@4݃x�C("��[6Ev�9?�����EE�PW���Ӓf.��pc��P)��'��3Pl�/A)�6�^5Ӝ �z��T[�}}LIq�R���4i��0�"�#c��*��I�i�+�F�1j~$�c�� v�|��5x��1��V���q28Z:�-ռ?]3F�8	V�0wr7}��Ȁv7����O+&���(�&�\X��.��˰o<�P�zq��r�`c��{�X83��~�K�B��b��~<��غm'�M����^tvw�\�c��x���A�φ��ɓ1m�Td2m�Aܹ}ֽ�Q�B�
G�֖��bJÆ�}{�zU�W/ctd�v���� R��9�H,��\,Y�Y�l�P�x����c��9���q�9KНՂ���]y�F�g�W�.@<ӎ:id�ě맣"��hd�LʟA?��۴E
c�d�T�Y#�?�l�j�ԁAu @��1u�Ċ;m����r��h_�Zn~^G�5�J�D���&g���vV~[���+b6��C�bD$���D,�F���mϺn�P�N��� ֌�,�H�eۧ��4I�	��a@=���x�G����GO��ҳp��b��n$]�M��>����"�j�v<���X��zl�6 </ՎX[b���sE�Ia`Q�"�3J�$����������~�(�v)����������'�:�Ɗ2i����4k�e�8'v�ء�#L�X�@�-�85�r�p�|>B��c��I��9h�5��_&�qpV
q���H�Ο<ɭ���KᔯY�Sؾ�;���{�v���z3����L�Y'���8s�E�N+��n�W��1?��-cx��w���U�7P�F�'�q/�ij��r�˨v9���?����5Z��.�X(}�t�Z[w���7��a�:�1����m8=�6���y�Ь}(�K���h�ƄM�uY�{���p|]�?1���ulY��i�tW�	3��}�9���25�JØ����8��#0cJ7�3i�<�F��n�PZf��(Vʕ�y�0x����&ԚID�ia�U�,�M7p�9��S���y}"�)���kw��G^��=�cYT)4�g�����|����*w�Κ��{�T��j8���~1��S:�J��D�Y����<��*0�P�+o�J]|3�B��ԉg�!n��@��t<���v1��7����L<���e3�uv�����˱���䨒��7APZ`L6)����(��kw��WNcꚵB��N*��Et�-�T�KO��t� S~o�p�.Eh���*���£Ϭ�L���,P*������݁�?\�&�&ѫ�-����0P�a��n�p��8�ȅ�>y&vw!���Z'#����6lف��l�K������eN�SH��K&�Ģ���=�b���7�_�k.9j?`zǣ��/���I�!d���":@ڬ�Ӟ�=�5s.F�6m݋������!d3̙={���֝��I��� '�r j���A�������F
sh�Q+�4��2"v��<W]v&.<�x̘>IH8�����׊��m�>,�mT�z�N�Z�#�����-9��Qd;'���Ki�o�6���!$bm�(���(��l6����J��vc޴6|�+�������M�m֕�1�r�x�嵨4����Q�2�E�E���r&_�IdB�x/D�`�=~�^bD��$������VK9Ԋ#H��8pf'��k�ƒ#f��`y�rӔ��J4�<�/?���x��5��(�8��^fRt�>a :�S+��_��`QQ��9v�9����(ǐ��o����៾|���0���^�+�[��e��?>��b�h�nzq���uT-˺Q����sr���7�Pʐ��z�m�j8;n�h�t
�D��h
Wd���	�e��*���r� S�����bT#�4�T(,��HP[&+�P����SNLUs����7�R��<�|I6C6��h���M���D�>պ��l�4��29�����#ð��j�BU��+��� O��?��I��z�H�PY�<B�A:+���{#�2��t����׿���~V����	�4A(N�R�bY<�Sd�$�i��y�ya��Q�E����P���"�r�	(H�jP�`�(��F!7�j��t2�x,�Ň/ĵ�\���@�-�b��7�n�������cJo7.9�T��QȲ�b�������%[���L�;�tf0Bz�<m���}��5�Z�31wU�	�?�H��:T?����+ϸ�:�1�/��tk�J���Nc��F�Rj�~KWP�֫��:�u�����CYal�/����#p�tϼ֡F7���O�Z(��=\��8�J$�iE�a��6Є�-M9F�y��n�shT���5sX4w.=�$�s���K��@#���@c�X��O=�:^~s=�o@�c��|")Ig��jˊ�L���Q#ثK����Z���j�A���p�Ϯ�c<𖎬]�	���`8(le�S2}<+Ү�~?���M���'�����$YL�:�)�6�u�_?�PnM9_{/�G��8WTwn�f�蜝�ҽ���DR��H�B��kes�[��^�����M�H/��(�H�,"�ajo��瞶���D;i����j4�wv�yV��+W�ß����Q���D��;摋^Oڌ���]�Yj�v��,����E54
�4vM����T�t�?������x�D�ckR�b�n�i�5�u���yw��V��_ޠ@���趞Lc� V+c@��5��
��8�[Md)��	��VE�T��Yf�l�\r"���TL�
DF��4v�p�� �� }���/��c�5b�,PF,^�oQ�    IDAT1��c	u��k�G��y�>�
�^����|��Q���c��VF�>k:��k�|e�h=�M���H���Dc���Ĕ�\�Le�`
I?Q���������xH�)�O���ܐ�l�Xet�i�q�F� o��,$��v��T�bL'��G:*q���#~�Z��2ǔ�e3F�Y*ך#�W�lp�
Le�jT��d��i��L�=�����<��s�ʛM�#g��]v�PyEc��z|�ǿ`�S����Wī!?���&.?�d\��L̚ڍl�7����1ds�x�`��vףx��U(5��tOF�"LAmT�yd�v�<�:�|���ڥG��_�ṿ�ӻ����D���)�g�R@*Vǹ'���>3&w ����U�~��xm�YTI��|\r�\�i�so��>!t�H�K�r,�ha����Q�7׺Є+��?�ȣ;��k�E$�UL����c�Y���3�����\���M�B�J�Bؾo O<�{GcX����n'�ǋ�V�H����D[:�J����2B�ND��%�B$혇��蓊ɩ.� 8]�U�Z�����)J��u��r�'�᲋O�Yg�iS'!��1*�bEH��Zvb�Ko��=����h�a�N���BQ�K�'����K �$�#%��.|���>�� �ۗlV�D̋,�P)��)�WG���9=��?}�-��� C�mOv�����!!;_���+xk� B�	x����a���	�BǤKEfz$G�ݭTR���"��S�/��-C�����Hu@&QG6V�Y'-�?���Bu�RL)�`��$��,0���0^yk#V�Z���l�{��J� �i�,7md�d�)�cg����)�@�XuZ��T���0un�H	�ēT^��	�>,8��|*/���Ն��tL5`�P�x&�(v�b!$�N!べ\Ų��ʛ��B�3/�#q�3��o>Ţ�k�TCs� q�Z_�8sh�J��l����5 �(�-2�O^s.N:j:�D�&WJsT!�!JN�z� %�?�$�6�րǞ݁_��I�i�,�O�V
hԊ��F�pF7}�������H�B/��V<�"FF��Lg�O�%5�:u��q�2�j�P��h�����vcd��T�G�i,Ƙ"m Ƣ��w��Xʡ�,#�!R��I�;kz{:Ĉn|l��Ø;g�&M@"I�Ɩm;1Z��y�p�a��^D)�{�����<��z��]�2�@����DL&�f�e�{N�]R'ЎU�@��q8
���tpDͻ�$�ϊt�o��������� �#�j�E�o�*���Ǖ�����v˟޹I�������{��K�b�f��B�y�Պ�^вD�ħ@D�����J��,E�#�W����b��"Ñ��&�!$�DJ*hִ(Ee	��c�×>{��F��~�+h�H1���B�7�a�p���ֻ�P�%�Ų�ĳ��Of�`�q*!�7i4���o�R���k�߉��ՔM^6�\��k��N+ȕ��^�����?%�BW�Z�9،m����rE�����-�X�N�2}w�ɿ�����p19~�č�y �hc)�#���S;�Dk�����%�~��*�FYg3��'gZ�▹���8��Q�u�p�I��sO�a��+��j�{��(k�MI�n����k�nî�<�>cI9'%ߛ�"Ѻ��-o�7F?V6A=���^��y�/[;7���PkՑ��Кbv���H=�o���l�:ٟ�&�cD����A��i$���8p�5a�2��ဩ�k��z��F˧K�0��IE&g�r5��WF�+��ל��]|<��ЊF]��
a��ut*��F
c� p���Wb�@Ɍ|J�5=�/�\q���A���I�	��G_؋��n4⽨zID$.F�{��bfo�1�7�D׀7����h��o�`*������\P�Ő�,ϘD*0��ϑU50��x	�jCd}�ǋҼ��(E?��Z#S��&��(zڳ®r��I�c6��1���T�bĞŞU2$3�Ry�M��ќ䘒��Ga:��σ���0uT^ߌK����&��W�ȸ�Z^\yi~���\�?OL��u�?n�?����Ӗ�G�>���8����u����P���;�G��D��gO�ǖ��sO=��+��W`�h5�v��̐��O/J���]�h2�/F�U
�l%˪̃�G���Ÿv�h��������Ŝ��%$�&��Ai}�|���q�A�>캼�>��_܋w6ߑl�K��W^0��vJ���+���?.��=�LV�J��އ�4��R��c��
���cp�K0�/�i�9�|v�Up�G��y��	�pZ���K�:7c��n��q���.�yo'�e]�3g�ᔓ���'���,�U`ӶA�����ak?b�,�ф��5N�M���vd�Z	���O���9�1c��L�lل�k�����h�L,�?�m);���.�ȕj��èGR�2Ǟx&�l��O���P^L��"�L��i}}H��(Wk�30�=E4<��ΩF�Q���/��PWA�/j�K(�G�+i�p��^�����/�EY��i��ѩl�_S�W�݅7���PM�Uk���E8�{���p��\�d�T�l7��6u�&�Δ�sK���I�RF�\B)7���A�%���?c	���kM������ ��$s\�ҏM�=#u<��x�w�w��\��P��D�ebڤK+M�H[M��Rp����:`*>،�ȥf�k�J�I��&��v(}��G�)sL���L�L��_���ӹSJaa��nC!1?"0}*�)��6`J�Wg�����e����p���p�\ ��Bg�������r�*5����y��j��n�����>0�l�F�ذi6l؁�qN�H%��5k"�͞��am��_�#O�&�4i����_U�z	����?����ü��gf6M�]�ܹ�9���4q���~���f�v���Ɗ��"�� ��똝}�fR��ʕ���݁Q���/�e��i�;�J�aV�V1::���0���g�.]��j��9$��d�s�eb�k<��=ԣݠ�Q$�fc|��-a�$S]�$�'����BȺv�K�b��a`ꦕ6�I:����K<��0Fl��2������MT����Tt[n��t`�L�7Ա����*
�+^�5��TSsni1�	�I�G4�q~�l�7�u��O)��UI��?�[�_�c�L:i�Vt��y���p�xjT
��I�4�fa�{S����q�Y�c������>��5O��{��i �wzx��+�쪵X�uP�jD�K�8eƮ�]�!�$�MM����615����,�	�2��9�\)h�i"��zNk��lw��E��3ѱ���:c-i���?���B��V��5�R���s�0P+]�=���/��;jc��y��"ӵ�a��"�f�%��H��˚d%�|&{����Wת��
2��*��H�B�1�G:g�v$ԍ	d#�~�r_�MP�%^1N�*`��^x�=���3�5\E%�F3цF��H�T,�N�-it��확�kfS�c���r�l���p�G�����5��q%��]K]��hw��D`���4��&�lp������;���:�4Z�c�7��-��lHП�7�U`�@���Q]�ej(�&F�q����lb���p��K0!���y9�Z�
w���V�s�~[?���x��$zm��I����p���c2�^4cF��@��k񇇞G=�(ɴ���~�](�D&����&W�����QF�Ɩ�6�`�$��Q���#4���<��ׅ��ӘzMчV��h2fO4�
L�jQ�����?��R�X0�G����Тm��+��{�ƽhߝ�&R15_�����(0��4�`ʈ>J�L�64�:#�W$�Nc�/�b9������ӫ�+�e'����p��L��ׁ_��8�{lB�4�����9��ڥ�IToꝏ�����w���ĉ���+8dN��v�,�٤�NN�Arŵv?,[Ϊ*q�%§���=�w7�e�6�Ғ%�������7�_$S71-5ø큵gSj&dr�H��y��g��W�q:%�T��=�?����w�"���L_������y"��ύ׀��%�������2�qsSM&W_�O:��<T���99��|��xd7R,����Ǟ�޽{���Cp�ዐ���Pϡ�M#6r�G�s���o�˞_�m;�ʜ��瞀�]�f��a���=����g^ע�z�d�L��7���]v��k�h��q��1��Ձv�ٕ����58t�lu�L��k�Wmċ墀[v=��2FK5�P�0}ޡx}�V<��s�EU̛�˗��E�E2A#-�mއ�y�"M+��1�Q�K!7>WX��夷���ם��IYt�EV/#7���<�d������U.���򪼻eO�z��!�[�+W�"����4�\| fϚ*[c�*v�+b�P�JTᣉ�DSh���{uɇjT�{!�drPd(}u�(���Й%���0�6�)m�IR�f�#E�ְn� V���lڍ�{%�'i�#�A"�D�XC�®Q�j��v�!�;O�]�X�!��-,%3�i!~	ŀ��Did�nNE`�lcRy�4�RZ��*u�3�O�C�--��F+�t%m��N���M<_�\.�Ҹ'D*oO���R�f�5ٌqasPaT��><.&H���7Tv����"P��U��q�+�#��4�zq�B?��
[8�� s����-�X���X�a7��
3�t��`��I��g��5��e����л�l|�M��7KHz9,���Ͽ�t�x�Z|��b��T�G�]�s����w���P��U����MND,���U]'i\Ap�mI>C���!Lė?s9�#]]'p�F7��B¢-�a+d������o�O���p'&�> �tF\��}d G�Q4�ԁRW�b�*����d�LN#�
o�0ц)� ��sw�N?(�,s�T'bOf�g��A��0$�y�&�??>@;;��u{�vέp5�����)�d�8�,$R"cQ�Z��[�k���D(�I�4��Ж�c����0
�d�t�S�z㏈���\�O˾e���92�Ȱ�s�(ѿ��x��#��e睂3N8D�a��j���>�s�X��y@�ϻ��Գo���WU��v��Y�E�u3�H#�6Z%OU3��i[�f�t�(cEo����p?*�]qJ���Mu]�I��S���h�)�N��dR���R+uN�:aUPh�O*[�z�����	�T�o�j����������B�Mʕ�jٷ�V3��ј�-����؈h�])���~̛=�y�h/��	LCc<�)3U!mT2h|�a�p�u�f<�b5�^�Å�8��1x�8�d���g!��	�Rsݪ���ۭn��|�4��ko��n_�L< m��ޥn�JֵĦ�{6�5Y�<?)�\�4��y��0�h'm�uqCRۈ�+�o���e�n�}�}*�[��0������`y=�6&�>d�Y��`�>���Kd⤎�;i!>��S0�[�<O�6k4s��P	�����pcoYl�ï�n��cy\~�y��0}R<]ci�ʄ�S􍻀��$^}w�,dC�PTn�G���؆�ϰՌ�>թ��I��C�Tk��rb SRy#�1�0ǝ�<��Ε������V��I���D���)=>,�L�ES͏��i��K�:mҬ�ڄ
�!͓$�TSi�c��I \��Ĵ<Zv�Ӱs�����j �/�z�	rM����A�zQd�m�.=i���2����1u��Ww=��~��i=�\��t��z��~������ә��f�W��������ZA���f��T����8!�`�׀����O}7֬ۍf�]�)���dBh�1�Л���\��/>
i��dbz�����?��z������3����O���툲��a�`���{���MHe�����*�⢓��kNA_�lS���c����+T�N�B�!�nƤ���ҷ��߃#L�׿�1̟���i X���xk�Z̛3��r":3$)�灧�|�ٵ��}_���<��U����e���k.�uW]��@��_�q~���Qn&���C���ϰ�١����a��霖N�V���Y�*G�3���7`Ӧ�8��c0}J��@T�>��UnH�����;�NO��/��S�^Da��T���KOƵW��)�zq�al���w���՛�y��`Wwqx�)����IT�#rj#�<�8i.:�8џ�cZd���J̝=�@�Z-�����%0e�b��
��e��c��X��u�Vw�|�sWa��y�bxwc���y��8��b��!�ؠ�� ��p��T���N=
�q���}���ݵo"�ᯮ���:}`*�I��Zs,T�ʤKoٍ���a��Q�~g6n@�RE�=����%G,���	ؾ�_��6oD3���$ɄL��,��V�����k�;��`�Ĕ`�O�CHO�s-�[+Sř��.��5PA^��L�h�$����(�u����i<��PDnpXrL	�#��u����iS�.�KpbJ}i��(jLG�b~��c���bR#�N4�CDW���K9Tr�Ȧ�>9�3O=�� =��������O��ww!N�;�)���?z*��d`�������ߐ�"5��PS����H�H!�E�I����
L �n�h�]��!�&��� �u�����{�=����O6��R���z0�W(:U��l˳��/-E�6�1�"�R��uG�M�>:�?�v倿��_`՛�Ќw�g�D�i�2q�05+n������D��H�-����Thp��=��u3
��Bg�D*]��i:��Ũ�����&���4���N��(8�3�S6D0M��~CqyWgYNI؜%K�Z΋���$ɤ'�X��pv����F,6-q���O(�����������x:��u��ֳ��}�}L����
�&�#j�2���:)��2==��#���p��vi:sm9	F �TOǳ�ӱ��ֻ#x����ӯb��Qi�&ڻaS6�DC��"�D� �f6� �3QM���-���ow.�����ܵr�e�a]!��h;�6W5�z�$nȞw�呲��:7�h��(����
l�{I��Ie�f_��驽�_0�mv�Ic�ϖ ͒e$jL��=�X'� ƣ*1��+�V�(���K�^�+#�U��q�Qq�9'b��f���o(sE���6)�t*V�u�G���W���w��b5*��j#�&�15�["�v��,��S���1��&��Vy��F��wפhٞmwr�K��\���4#��Uc
i&*^%�J�F�5���r��
�����s�<�&��[�}��sm�IN�Ͽ~�*��K��.�}=�<q~�߳󗱑�qz�"��"�=���e'c�����F� \cQ��[� �]r,�v}�;��Bx��0�������[6�l{�=e���?���������Ө5w�{��/�gR	��m�O�����w[�ָtϬ��	LՕ��h��T�va��Ĵ�������e����*"iRq��HFш�<o�J��vMjDc��h*��>jL�"���kn&�XW���F�(�����+9��
���P-
0��f��]�n"!T���#71U�8��kV(`�����K\�ӥ�HK��0-z�G��_��n��S�bi��%q�9��.�g:����W����U�#aL��o��\}�I�85�
��X����-W��1f�mQ����������~r�nF3���͛�P#���&����q�EK�b�?��q�o��?��F
�#a$u,<�����p�̤���!<�l~���0����K%�??�d�������ګ\�u��������djJ��l������e��{q�	�_����yI�d�W��W^CWW'�9�4̛ѧ�w�غo�5�)뷎�7�O=�2v�B�Ӧl������IC��é?�y%~��O    IDATq˃Bo�4=��gv�N�����Y��F�#��Q�M��
���	��V��-��ಋ�G�]
˖UK������Z��"ظ�k���H%�W��o�'���>������c�%�*���}u��Oc��[Q��]���4m���Ⱥ�tu�n)��v_��"�w�\�E�B�۱y���p�|�n��-<�����ۻ����"��lݲ	��.��|鯯@7�����s��/b�s�P�'��L'Kp��alt�0�JJ���7^�%;�Jި �{���[o�C¼�3�<�6���i��!�o��g_|�mهW�l��]�����Ø�T�p�8��>������ӛ�{��h)/��&5��\��,��G���Q�˶c1@��=Z�Rg�i�PG-�TձP����R��hkW`�͠�Ds������]7���3�(�H\�)5�O�u��g�A�d�<:JH1,��%4��ʫS�O� S���GH�f��a��Fy��p��Y��W��Y���+��v�7�/�s/mD*����m���Sp�)=��g!�o���Ux���(63�y	� �#a���+#\�!�R��������}h���/������7x[��䁻|��mR�ɲ�ʄ�fV�\�5��Z-�Ji�?_���D�&�:_~Hs�2I��u�}��>ÔЕw���oބ;� ���>��4,��6��8��ЉN��_W@�+�LE�^�c���(�`7�(�-ӭ (�p��N|4gE�NY�?Jv&cj��:1���.r�Q�I��կ�):%~��h#�ŇL��06���lĺ�C�G;Ј�eFD$��W��rSl�}|ஷ֟ˏ˳�մ� N@�� 9*�	���� 57�T�d5��q�6�^�*�l4��m�QC��G�Y����Im����p��aBY���FX���ZJ�T�O�<�6l-`�ʷ�|�ؾ{���64��
�`�0)��B���	;���w����S��̌��~�Q�w,i(��������kj؛(3�+��[�c���/l��3!���SXSƭm��>�?�f��5�����#��?_�������4:O����'�(i�\̄oVKȏ��QE2R�������ca�A}��К��`��8ʲ3�a��yg+V�O����Ј"�hC��80���pT����\�Z���%)��~��0 ���u��`0�����F�!k6)K˨��3���Έ���Sʡ���(1��k�Y�x;Bє�}�"�N45�	���k��+Ly��6�ϹxA��׺�-ʦ�.>J�&���g��^����I3�4#����8��ni�J̚{=;�F=���F<��l߹�rY�Hsf����bɢ�1�/#S�HHY2Mf���4��ks�D���!e=�����s�;F�K"ʸ6�M�CɈ�6Jl����d�{+@/�s�U��k��w����u�NL[�i�C͇L����)5��Z�͋���21e��O����e�H:;�"�?$T`z7Ĳ��R�Cݙ'��ݖ���x���LLsC(���&G2k����cڐ��L�9����&��@����az)0Չ��}�Ӫ1uN�-�������M��{��=!�xo{
W�}�Yz�����z����܊�xM@��K��~�8d^��}�̱M���U��r>�A7[�1�H���l����{V�ֻ�Ů��8�rcK���;�����앸�%H�LL���Mw��P&�/�D��Ew���E:-)��}������^�7|
K/X"��G�\���|���R̛Շ8MY�|���P.�R=��V��F}�F��<��~�E`z���31��Y<�^[�/���,�c�^������kF�󭋜�����i� �?�Ϯ\���q��QdR|�Wຫ.�K������'���cud�'�o�l�S������-pQ���#���^�g��2�M�ج��ʾ\��j�����ܔ�BH#�	�{�&�("E� bEETD@E�� @�%�@@BB
�	���g����k�=3�����<O$&�ޙ9g��׻�[\ޚ���ކ��y*�¦���iڀҢ�c�PĂ���m�J��`�Jl��	o���!\��sp����e
J���6���%,\�.h(DWQ��ִ6&&��Ȇ��)�櫾���oEX@��lڼ�>ۂ�3f ����訌�� v�_���]���9ذ�Gbb���Ku�着+�s�����L=�O���RT&�H�H �|Y��(�0e\=~���`��	ur-���1w�\��m��wZ�٩Nz�9�~���M[z�����MX��]C%�#���7|�|�m!��;8�|S	w��6�ȣ�ݗ�
b/-�Dd�Qd(2<�Ę���E�k:�|�IOᆯ�4$���k[�>��)��E��C��B��ub�GQ��s�T�$9��^�t�����b]΍6X��q1��3҈�����Ii���lA~���i�P�U������G� N�n�^�?�х8���E��_~�n}�|��31n���Y'���:A�1����7�г�`Ѫ�U�H:'�tr.����-~����0�I)OZ~�W�,e��"�]��u[�'�}����p�hĹ��!�J�̬f�G>���	c�p�w����n�%�}�jKa)M�ajy/GS+����݊���$rH�� �a)���T�^Q�������7�Ě�j�S�h]5J5MR�D�躌ɘN	k��1;5�S'���3���U�$�@��:)m����*a�A����-\�<��v���:�#3��R�w3C�(�7\�}'�ŉ���k�}���*��	`D�/�6��:l���d�8a�z�f��5�^zM�Z��Zd��/��5S�ڼn��٬-�nQ�<=%N�r(S(��p�!{�S�¾S�"�u'�!�IKE׷y=+�I�gۀ�����l@�D9C��b�g�����?�/�ʐі��<3-xW��/�b *=)Y�
v+��ҷ��*��<�Oa�p>�u�TK�Pm��O��ӟn3tuQ[)ծkܬ�]־�z���iCU=�lF�Nͪ����T�̘4#�
yɏw����Ө�����K3�w�>l�5��	�~&��R�b�{���C֊�}��U�����r�N噧�F'��A��3��)Ԝd���dʬq�?�e�^/�dbjB����SU* ��k�b]��3��c�����*�E친��&��B�Z��1zd��|���6m�E��5\��ۻ�vaهY��JC�L�펧�E;]�^�Zɓu �ZÊ�j�5�X�bܧK�I��f�)�����q�%�b�Q^I� ����3����)<��;x��y���H,�E�y	��8��i����䑂?��JA�Lr0 �����s�cxe�*<��"l���nυ@H�7d/3L����3�z��j��諍9��5�T���B/����`�i4"�h9�ަq%gj���χz�_9E��:�
���|�(�MML>y���4I���k\�1?��`�Z5\��*M�^�t�F�3��x0(�G�|A&�ف4�����	������0ƣ��@�ɐ�J��Ԙ��}���cj��W�7`�_���2�����^G�9�uQ�w�RyebZxb>�xϿ�I;�=��3�K�E���k&Ϩ-�����v��j�)f��-��$8]�1�;�>o�g7 �)�C�L��F����ω��Nd�<��*����0�� �05�۳w��J�;6,"���!����hk��i���=�����;�l�'�o�$L�<^6G���[��џ�a0��,nH�B�H>�l��tN;z~v�w��0�Sv� �Y�/[!���--c����fs�f�U$7��v��0�)b��,�d56l�&��X�/���Gc\K8�Ht�>�w��$�]$�Faب1F��J}�:����јӀۏI�=���1~�R]׃t����}�>]����e1m�����G���O�� d�u�`����ғ�`ރ�+ע��S�F4�q�5��	G쇨�^��Ú�9�������.�î`�(������, 2AoM1�^�5��{��fSj���믿����{L�$���[���JՎ�PP}�8������'�b��D"dR��v��O�/=ɰnLEO =Y������]��p#�A���^��A0u~w�e�0��JG�}~�����!3�!V�SM��=4�n![ ��d�|�c��ҋu[�0�q$�3�/��C�­W}#�}�0�xО~y�l,Z�Ǔ{t-Z	�ȋɟq���m�R���ZT*�P�H�ɸ8ũ��R҅�"�(�u<2��[�{ ��}b�Jđ�o����2g'�v���*� �m*�Lw/�NLKj��� ?���[.��A��y]�~�����ꇗ.sF�D
��i� 5�R����1Pn�CrL��J�JjǏ+�/���O��>���&yl�	GL��]t2FRSc��}%��7��_�` RC5@��=�x�P��!����ӏ���cDS�hH���֨�n��a��M�x�H�Ig��՗��m�h�l�ч`0��L>�L,z-v��ȗ�5@
8��=q���1��	����lњKi\�V2�^�Xsr?��l��S/���� �&����СL&�f��G?��R���3,���~M�^�嶅WU�푂Ih�5:�:�Ti�����p�G��*]���_T�F�i��6c5�L�D* J�_tU&r���H��V��<�ǊyZ�k��m磕%��� ^���<�6�̠�SWv����c+|/�FF�SN>�Դ�)��y#��`u�R���q*��&����4K�Sl�j� ָ��M�g�I���]Yu�'U���Sэ8��}q��a��i�cIK��r�u2�D�y$œknGG�/^���âO7��//.��PR��Hgc�Nqdf��(ǰ��lQ[�+}S/�L��\7�������5�{1T�vro�/���(j�X}a�����|��[�U����l�֖�1�7晵��0
���p�@4���:5s��!��R��#��CȦS��T{�3<����}��}��Ǹ�4$)�0�m{4�Ir����t ,\��.\���6`{wpe�Gĸ���z���Y��v�	v��R{4*�f{W��.����QI��U+	���<��{��ͳK�'Ȓ�P( ,�%^�q�L�Q�����ǥ�������<��4��?IS -�����=Jp���Z��4��r�3\{�+u{�ڒ�a�������[��Dݯ)�b���e&���+v�#8%;c ����ۼ�ۺ\��гx�ݥȖʻҨ��a<�[H�\B<T�ч.� S�7	�Gj�ǔ�'��6d=@G?�k����s��|e_Xd#��%��DI��	UYWxU�mM�t��cBdA5tga}i���D�8�� L9�$($��!`�BY�4�::�K�ʛL�Qd�PЉic<���<�b �s=	L�q�@G'�:zQ�$�7\W� iL52F 麈|WÉ頸�f�V��4�c9D@��f�Q�)�!�'
KF�|eO��!��`��ˉ��x�Yh�oT^jL�?��3������1�>�sO���O?1v�K��g�����T�����mW����t󫉚f�T{٪HD������+oWOx��x䙹�l{?
3]x
�ĵ�?_=� ����� <��j�u�SL��Ε�[�����D;y�Ĩ�4���`Z�D��~�b�|A&�^|���`]��?���A��K�H���r�ê038���.�w��C'��7]��c2�#������h�R/���z���׋L6��PF��Oh���1$�u��o�����՘�`!zS)��^���{����N�L��i���1m�*��T�y�j��БV�Ϥ����b�p���M�}d57q`0����/̟�.��A;f$���l:�r�҂��x�u\���ޗF� ]�a[[/�;z��2�%����'��>Ҽ<�ÇU[r������v�=J���#ҍ�T*X��s�4����<F֗q�5��=��A6<�W��/�&�Gu(�H��f�6����FF{w�̙���nEGO�C�f��zp�g�����DX�'����~�l��4@
 ��摡��P/ʅA8m�x��v	�o�=X�h���q��G#α�aTk[P���ޓ���W��O?�����5���A]ڴ�pܡ{㶫���zڧ�P��Е~u�l��h\_��R�����
�ɉ���"�R�c����6@Y6V��21����n�%�WC�]�b� �~ʑE��_2&eA:m������A����T����i���l�`��i��5+0B�u!� ���
0��l@���k��β�HKℇYl�<���q�1Sp�5�������?�-�*Tk��h��ԉ��������G�Ԕoe���m���*�%ҳBrHЍ���<�N
��N�%$"����m��2\O{ͤ�``�~xO!��,�Je���z�S�Hf�ȼ?�̙�K����+�q��", �!�^�r�5*cz��:�;��p�U�� �re�]l�Ķ�J�|�8���4�X4�tQ�������N�l��_, ,�F�'%��BUh�քH�^�	SY�S͖�j��^�pɴO�������&SPy�l�R̈́Ңg3��VT�����Ď�>'7Ӈc�?�t�Р��������X�{���}^x"��R_��q#Av:�j��b�R�S��T�xM����k����ΰ�gϤZ�9����RK/P�w�U���2�CGJ�)�<9�l�×O8��|�{��^;����zE-�añ�ذ=�w�ļ�cGg
�<�Y^��H��$�v�~Y�
X�����{*#�LmC���/P�s��SQ�� �Y�Ym�6�,K��A���f�����~�N��-�L�Dk)���+�*R5� 5�S�4#�t?��_����W���ԑ�j�z`W����J9�hڒՎ��9�ǌ���ӧ��}v��Q	��FÆ���Y}�f�(���ʠ�t��!�aэ��n����r�R�üf��sQ��N����������6�,����V ����H��&���hs�0*�Z�R�(֋|!'�F>������.9��|�d��t��d,2����+��k+E�ɛ7��Tye�)\}O��V9�j����}��fw1�fV���P�r�WUB�+N�X[��)1�`�_>jn��d�2�[�4T*��[��{f�/��a�)#���S�@7הd���,B�4.��t\z�i`��I�4ªՊ�}6����;����bsG�H#�a�����&X��U���1`����X�/τ����hK��h��$��_ T_0r��^|f��7zU6�ubB�)�+o�?%53������!�Ɣ�#}�t���1-��߮�G9:���`ZďCrL���NL>��@/W�sL��`�A'���(0Օ�=�MZ�>�g7)��eb���D�<�����GԎ�7�,L����:1��Y����q4����{~�=�8ry�3��f�3�[�T
�k�TՃ��� ��O�9x��yxu�
���H�AL�/=g��"�]�Tc�U�뾧���DcJ�o(X�n�b��sp���d�ÿ�ȼ���	�N��.���O9O�
��%ǟ�T(��^�w�0�'>���rL��v�;:��e��B�H�����%g�)8r�#ѨĨ�&I$��bZ���-���,X��B_9�X\���0��d�`z�̏��>���2b��4z4|�h�@x��-9�NJ��_�ä�1q�����ןƿx}��ZG���Nr���n07Q�7H)e>��Jw��%k�ڛ$�fTK7_�ľHr�%4H>٘���{	�n|Qq���h2���:�]>�gۈ7��M>�캯a�)��I����P*�9/��L6�#�8#�7#aA�E�n��XdG�=i�5	V��@{o��m�ζm�����%_A��h"�p��T    IDAT�ʒ��!���r��LQ���Ẍ��)z�Џ��+�t�0�l~��ذn��>��g_��8'z���h�Ã4�+`p0�M[��3��L����o���Uџ@��	G�ۯ���t��) �����`+J~���ʔ����3�[x}NlN�)�=����E���!�5���ܥ>�O�)'���2 �H"1�	�D�fbj�LMZ��^��P�d���F!�I^I(1L��(}���J0m�Ys��0%����7_�P�8�e����S(n&>�O����83�Rj.;�0\y��H�0�0^zc)�|�llۙ�=n,�Gc�7\u�=��<03`����` ��㓌d�0v�i�F�zf�W��lp�Aۄ�Q�6Z,p"�S-��kʼ@���A�#���e��%���!�J3����])��P*R��H���{2�}=�h�!$
��I������%Ac`B��Bb��0{5&{,Y�Q
�]:��T�/��U˄4�T�"�l0��� �iqQf"c�p��RH��gkx~�%)�-UI]3�T�_8ԔZ����O�+�[�.�(�H��{ �Pi ?�}�'��_~�(��Y6syΙ�w�c6wQ
�����{
'42� b&��-�l����������D̂�J��Ųװ<�铝K��q�5��R���+rQ�����ʰ�kr���1�T_��,Z#8��Cp�Q�1i\��l��Vl0P_r�M��0�(� H}k�*�6wV�ކ�iqtl�����C
��eeA�� bS����&y�1���<����er�T��6�H��͖���
��Muiո�FT����`mtH�0�P�m#��9?�Y�F�l��1db��F3�������=��(dH�t�q�������G"�È���gw�8`2�<t_�j���4t}U���<\ �6o�;,���,�8���	�#҈г9�����R�f������ 3)�h��<���k�ê�S�}Tv��υid�5`�0�5�W�>�SJ5�׃bv �r
{�K�o}'�N�(�9�}8^H��g-ì�!S���@L-�7�Mߓ}���kv�j݁m���5����T3�[��L�`e	�}��E�©)yI�Eq�R'�>~?�t����Y�y*�e�����G���S��?�����_ʥеc3���bA�w|����[��GF4mo�p���T_���>�6w�P7���ā��u�4ɤ)_��V��
�`_�ee�U��9��*&��L��y�pjʯc\��2ԋ<S,j�!l�%�~�1���Ĵ���`6E���o�G9�����v�ዖxќL ��o�@���L^�|�P%���W	m���Wv���4A9K�^d2�(��7�W2XI�-��:�<�Ƭ�q��G�CU�Θ���陇O�����jL�_��ϼ���_�K�iCL����%`.KS�fぇ�
����?�z�%|�ֵ�NF������/��]�F��$g�� �[�O��6m��`O|�&����9[  �X��Ӈf��_��2Ny׋`$$#%�}�����#1�N)u|g���ڮ��/�1cr�W�m�Ss��F��dI%�����:E�b�ߍ��6�����'��.�đ1��y./~�4H�$F��Tɛ��b��
R��ax�����Y/ag{;N?�H\��1�N�?c�������1�� �0�Ǝ�����@>���ص��<��Lj���_�GP��9G���>�=]��ڊ��:���#�� ]�VG�pr"�HS���Z����o���#ඛ��S�; q#V�[�!�;��t ވ�8���=��:P�˖�0��������`j��eb�ܜW��u�1G�.Gĸ���m�`m6x{��܅}��,��+HǕ�W]��E��F���,��c����	0��i4C2I�)=ݝȦ�ds�Y��o���*�g��]ݝ;۰����'�E��Xp��	L��Ђɲ�\���%��֣�	cᲵ�D�j�zd�=8������EkM��9�o�4���$�]~^� u8����j��8�1-�L5K�2��)�c�`�Q7�E�tR������y��@*o����A���d�M��J�0x-05�^���Ԙv!/�ٮPy	L%�J��d��i�����t��N�dZ*�~f3=2�f5���TR�!�'׎���n���21�Ge���܏�;��m;�1��(%�뢡.���.����1��20���럯	0u�ttf�W�EJڼ�QA)�@���y�����?��O�]�W��%iK^�����vJ�.bb@�S9�A�^�@0�{긎��EA��l��Ԥ2I�3�����\IO�m���0{�A�^H'7ٜ��6���V�M�hi�vf���c2�1.ʊg�F�Ƅ�j))�d=>�DV�O	S@�����t`k-�����T^{k~���d��-�\��Zr}WrOhV'���3-������˱�:[�|F^���K���'���u�׷"o���_�����A�g�L�����a��F7U52E�Zxjgr%�E��TWk��^��2Y�b�\�)�jO�a�:<:��|�Q�TH#7�o�SǷ�䣧���0u�4%�`G�T�Yu��קd�Hý���%�w�O�a����֍�O$	��4u|l��n/�A6���{���f�/.=���`�N��_��F*���>�a�Y�fro��֌�9K��	��;E6��)�i'n��p�P~pXf�P3�۬�,,�4�M����&g��ˠ�'(- �h-T�,�q������~{O��S����Qk i�>4&>�R(+�aWo	��m��O7aѲu�ҖB_�n�t�PX3��/��R��8���^�L	�,`mUU���:ޅ	�aIz��k��J�F�Ij�4;M�i�$qᦄ�Ԍ�l�B�� ��4߿�T��pi~k����^0�wŖ2���+X���r�PD'�r�Vahe4T��ҝ�xk��N�E�m!��\�����<׍����h��5�{��<�-g ��N|�����&�TB�D�%����
f��D�\n0�Ĉ���yJ-�Ӿ~��D؏�������-?�^�	��?���r����~��簡-�t)���?L�Ґ$'�i�e���3����3���6kZ�٢n�U`�1T޲ R2�ј�L�ҡ՟'P`t\��TF4���H��LL�1-��l��t�-
0m��]��\�Ӑ �@c�Pyو�U=��,(Q����l=�f�H����L5�OdI�<;*ِf�H�T�Q�o�����Ĕ���͕���?3�<�*\-�	�y���̣dbJ:̟��y|� �o�&n���3T�j���ʭ�:C��ʗ��X˶����,���,b���h�&t������Q\y��8���+�lك�Y�{zQ���8��-��a�)#qɹ�a��"��/ғEA���ǚ�*3����[�xy�|�r3|�:$�6��Q͞2S��P�ڶ"߿g�n��B�k
����Vh+J��:�U���f#�׃L	o��c�c���8������/Ds�G/J��x�|�M�J$��BCk�vj�r��8D�FC�T��fz0e��廘0�T^�8�8T�S'h-�*�$�=�|*�]����^,^ه��� >^�u!�⧗�ƔS��MWl��y��w����<�H�N)snY&�(e�s��[K �����wr���{���l�6��[�%�b�e�7ls�ż��K��5xj�[�����z���o��|E��:1U`��Gޓ�i���� �#Y��yww;2�xJC8�	�����p6F*�5�����OW���B�	�s��@�u���ЇG�}o/��D����/Ǩ�H���/��������ż������v��:��6��y�NM�F��'���4?b�)͏,��Zp�ab��Ԙ��h D����i<,�ϟ�v��r*P��J!�Ӌ|:e4���֙�n�v�f4����Py{��-��J�@���LL�d:�~y/������qФ$�����-��[���'�wI�ً��yf��F�h�!�����Z�5	b��[p�Cs1����B(�=QX��k�1��JSҧu�f���&�\J!��fLg�t�X��}������5$4�\B���#ܐ��h�&!�Ѕ@�"���`p���;��St���]�E!�G!�G���s6]d�k�Ӧ��;) �ȯ�+��1�=N�56�M��UWsd��2/S����	d����4`̩#/Y5�)fb��R����ފ��}V��/�Y�I��	��q�B�K�jTR�}��,���C)?�:� n�����������@΀b�9 ��E+�q�����.8�a@�NQfi�44����2+04��mq[�[~deNi�F$�s��wz����V��%5�Л�T^�E��� [�\�1S��ɥ��<"?�`)�1������q�9�`�--B��{�I��θ������)im��㠣g ��z�f�,]�?�@ߠ#�w���<e�nP]'��"��rָ#��a���7�H��J���t�յT-��*
c���<.MΕu=V��:���إIc�yk�������T�I��8��Ҥ�q�-�:H^=�d}�m/!�)�)1-�<�{L����1��Úb�4� �5����T�Q\�u+V�W`٪͢��鴛����/�r�(� 3E��R�,��Zr����]���);1��t�f�~�1Ū|uM�f��+{E��`u/V&��\&'C��^��!�G3��8j�($ث3zn�.����6s1�{})����Q�dĘЭw��w]Gjg?��ڊ	��^{{�O�i�^:X�#g�.�T܂��U$dq�˦P.�v�C`z�iE���fqz1Xn��\<��"xM�D��G(B$�i[z��� ��b�{+ܣ���
�{T�}��W@��5<��{x��M�{���}�OC82��>Q(��m���;�L��QѐW�E��Ѯ#���L0�!i���)؂�
LuIx{�{*�Uy�Py�^1?"0��4;���[&����(�X�9�28�ae�%D�^јrb:��)SS6�Bu����]�{����,E���*0%X��T^�(��ŉ)�f�U&�	����q�1�����2.��t�eG������ϼ&�tXcgs �~�Q������{����_�����:�$��a��]֞�Z���k��>v����I�vF����[����@!�	������؃�
=�?����Y�qσ/��ĄK��S�����qڑ������Ð�;X�h%/_��TɺzL�8�cF�ik[�n؎�k����(V�t4Rm�Q$�j
�$$�c�&d{���Sg�G��Qq��4���g6q%�N|���t��^i��+%�TX�z+��>�,��v .��|4ŵ;ǎn	�����g�A�_/�41b8��%W��DS
��-��ez0�%�?��b�ccE��J�޵�`
)CU�Udo���2W�a����q̝�4�Gpˍ�ģ@"�Ŵ�n��3X��E�~X5����ghz��|nN���(n��B�5���bU�煢+@\�{��n↨�����͉�K-g	O?�~����J� ����*�a��;���w�����w�����Q.��Վ�P$����oK�����LAVy ���Tqz1�#��u#e�Oh����������_Aw�Nw�t�z�e�D*�v���/����]���fb	0����T�,��T�VS)���A������Y����`S��T�8J���rb��Ĵ�O�O,�9�&�Tu��j����S�����ðgڧ3ǔT^�T��ЍG�,�9�+���(T��^�J\�vUs�(��R��fs-�Q����߇��FLi�}H�ȥ����8v�>�Ԅ�9f�m�kk�'�C�����8H�I��J�U�/`�6��8��a�|x��H5�(߷jg̺*�������Z�GE�i��ˤ�"�A���*�zt
���M��y�@>E��,1T�98pXԊ�?�:V�j9p]٧�J��u�)I@lס�F���uaD�muʂSr0�� }3���U�ZC�4���4.-u���P�`&����2h��V�b�?-�M�	?�L�M��F�PS��Nd�qf��R1���d;0cb�^��;�^��:����)6hR%`�N6����+����� ��}9晖3�(�j���<3'2�T��j�+��*�Q��(�KT��f����Ԙ�	�>a�9��~��5�jCZ3��(��`/��A�6G��Ա8��0�=��f%�#�iX՞g�`���=�L��ƨ������۱v�6�\�	��v` ���"[n^2NH����F��	2���a�f@h��NY����ј��Zq	7m�D�X3���YU�g[wi��v[e]�Psm����"� ��:E��	��[ɢ!]7+�ܸ�!ZG6b��1�:q&�֊�F6c�0?����i�y�q5XD����mdb��Y�n|��xiP���yQ�p����K���� P���be�l��,��G��mx���N��Yޕ�Z�ij���b���Ġ
���|�I�6�<% �NK̓�퇯Џ{���+�Ì��%��!x�iVY{��[kp��y�d�M���*���L���i��l*�/ S�\�ud]��K��l�C�-6)�>r�<��@`�t��S����N�J��bpx�����>� 9'��?�dKF��P���'�Aw��F�mǌi#񋛿��ƇE�%#��9P���xK�t#�m@��ai��n-�uʬM������T��g������He�j�9+a3��'��
0*o(���'0�:}�2,�7X,#�3��PZXG����Q����)R���'�/F81M���f��P���(�@"�PS��t(ѡ|�(@ڠ���LL�1�k�*1�c�0'���r��;E��њ�� F��ͨגlA2V��M��(�Ը���j����*0����Rc���Y���u����;��� S>�7\u.<�H�«݁Bծ��"�H�Q�򛯮�O�)�I�
 ���m��|�����d0iL�\q��Ҹ
0͔i���=�/ǩ�,!�u0�9�c��c��	��АL � O��>��>�ыt�E8FCS3�������PV6���.�aY��j	DC�CC�E#�KD�)�Ѿm#
}[q��ઋN�8����J^]���ұ�`�V;���3J�~���_�����g�\~�Py��B������b��%�>�4����`�G�i��(���i'ʛ�Ğ-��Ӌ16	D+���ת��|��(x���i�K�� o�G��뽏��Ec��z�r�wp�qӑ)�� /Vn���?>��{Đ�� ��t�����>Pt�,�p�0eL?���6�Q6u�"Ճ��<|5�ٖ�U�^{�}|��������>X��o�==;���}�_}1�g�k-���w����Z�P4*�^�g}�]Ȧz��q���͏����*]��<�Ԉ�R��M��i�M����<�� �^Y��]�;p�IG�ƫ.FKCP��d��_���ys-_�1�y�UѓPpM�-�\�j�^�lc��.:�d��.�7�ή�[�hN�Y2x$��甄ʛ�#���4�����!5��L����� :q�#u�ή�4r����������9Ȏ�9p�[���3K���"�Sa:мI����I'��d&�����=�Z͍8? _�'1��w����h]j?����Ms֠���e��ד�c��<J�$�Z��A
H������$���X��6�j�R��0`!+�6��=�
L�qd�	�3eG:�A6��>�˜��(&"fM���He]��T��s��y��P��=ϯ��@9�.�t����R�8��,ѶY�����DH&SF�a�2_�^X�*�0R*TI�Z��g����-� �k(U34?ӈ��Ry�Բ	du�ki���i5���ihNJ�x��^�9��3��D��N��)�ß�����򯟂C�+L���    IDAT�a�Y�9�sJ(me�m �Ǔ���ѓ��n��C�UK�7�}B�54�Z���:)d����[�6��L�Hdla^mH0Fe��)C�7--���=�N`��	xI�����;\c���B������� e��#q�3p��{`�	c�:<*4R��v��JE������پW���Jꊺ���OV�òU��ٶ���Ggw
9�
<;��dȪ	�F�(�W��2nb5,h�fC�=�hū�F�%�f�����L�h#�7�,��Z��l���0V�'����_��EAH�hu4ׇ1fT&O�}�����GaXcuq1D7]Y�f^5S��M@��Y^mk���՛1o�,\�
�Cy���'�2�@$!�_��Nj����|�'�SW�}J�Ǧ��g���ؚK�j�)#�P�^\m��!�J!,k��h���tJ�z��i�Ϻ�^�� �߇\B�~�?����w���1�yNZv�S�������_ϡc(_��@L"@�`ZK+��bժ�ea�T9$��TeU��iVq/�t^����D�Fc(.��]˺R�$��L]Ry�v�w��L�iHeb|:7�n��o���A	u�G���B�)k�#B ��`��.����kb�p��p�T:��McC�g�ǿ_�S/|��l�PJ���A�a:��sI�X��	�]I4��	,U�5�80���)Z��%��g,�*�6�J��L'��jTDG[�*:1%�&Ӫ:�$0UW�B�����[b�%25��	��T��:d�	T4�Cs]�RY4�Y澋+�SS�RS�f��W��:�29�ut���4k
�c�E�:^2�H��	7Ӹϙ�q\�VV)]�$.��x�g67^v���ҕ7MW�Y���so��F4'�����<�L���/Jas�㲯���.�Q�q��0�}��-
 0@Ͽy�^ƈ �E�w����w�y���!L��W~]�)�F���}����Ca���uq/�;dO\|�q�}�No�.�e�5Cxp����ZtP$�ii �m\k��C(}�ǯp�cQDٚu����ʩ6|�C�O����'K_>���.�`YQ�	W�m�P��H�6��ŋ����}��K�����Oo�Z�K��U~~�[x��Q4 �Ҋ�&�jdt�dw��i>��Nz �\�6�q�O/�8���1��ӢI�!�ZTg��E�*t���������mm3����8��c��D��^ĭw>��k:�Bxq�\�Z$)8���ĵ�_��ۮ���o"]+�(y{��YY�����G�L�q��9]V�S��o~�[o��zw�G?��\�m4$~�1,�i���g^�D�b�C$G,ӎaj }�(p���۟\(T^Qq���
��z;(������m���Ju >�&����:q�	��'�_���Qy2H���]/��7עhF$�Wi���H���Z[#IӁ6^���F
'����rb�.�k]#��@�)�E<L��Ӳh#��g��Ubn�pF���M�)]y{z�O���O*/�1�����ꈇ��y�+���B�g��4��G"�79fv��I�R=��]!-�l���;Z��سE�H{o�vo�︦ؠ�����u���{X�u ��0�-<����4�)�dRk2�R�����TCPmZ���{���UV\h���X�rI&�lQ���ݘ������2l�����}�Ҥ�A)[`��9	y�,��Q�kM3Ơ���6f��m�I���@*��q�ßo��Zp*��)�x�{�E�z9�I���F�hS{F�T�N�L�F&�U���Uڠ�Y�Ui�V�F�M�*��
k_��s�Z>'�b���vK��o���,rU��}��\�)��=�ӯ~���Z�ΔE�K��7H�@��67Zֳ��*�Lz8����]�������u��D���TO~=SL�G��Z�:`���i$�(:G$1������G y4%�2~$f��t�ޘ2q��I;��T����wf׮y�V�(�f��uG
?ۉM����mX�q+�;����/��PZ�u���h$��V+Km�X��Z�9�U�>�����y!�I��J��A�,��Ya2��^��(��X4�#���:�w��SvÔ�[�:���^��k�:"W����ʚUYH�ડ�r�ŉ��-=�ϢX�t-Vn؁�TQ���R��^qJf�eִeU��ґ-ؒub�`f֩�K��� k��6k�N��T��y�x����ᐂ<���=��,�,�A(TH�4l�eQN�#���K{����u
�<x��o���&�L�=�P�>k�Yoc��o��Պ����U����
C�R���Ul�weG�4ê5���T&�愳 ^>#��̐�S6R%*/3�rqP���N�n��$#Ԙr�R
D���x�u�ʤ�&av�ߧ�/���l:��=8`�V���HD KH�<%7�tp�O�,܌�D9X����	cN�Q�.��$�d���{5�|s讃�ʲ���\�4�3��l�v%���� ��o4"��d��V��� �����DB���SY�S�5Ջ��	�J˘!�L�����AK}�1?�DF�i^�b�������W&��2��O�s	LC���(���K}�,F�?J���&��Zo(�w�끅?sLU+AS%qcϧpSH�}8��=Dc�LF�3?"0����ҕw��F|���8�ˇK�E����f� ��sN?	�]{Ȱ��ț����.����i�x���T�}E������/c���𕲘4:�~�s�8�2�;/���z�d]v%�27��g�sN�����ʮ������ߊ�xw�#RW'�R�t�ڊ+����E4�W��������l6�B�έ��p��3p�%g�)`h���t�r1���Eg](�UD*�4!F�D�R\��M����]��h�r�%v���7�=7_wZ�%eqI�N�������P5"9|4��Mp��G��q�۸���K�A�{����[/Ǹ$)�&��1:yvXI�e�y2M�Ԙr�q���z��38����d�ek;�|�]�]�AhA��!��W7��3O@]LR��;\���'���EP;	L�;��],ʤ��(;)	n�s�:������&y�����A6�`(�C,� M)94��r�lf�1��L
�V��t�V<���x�����p�u���k.E�F�ߛ�}p>���EO��1Fc1$��S�׋��6��}8��p�O.xqA��H���ohE�
[��@��&H�U=�ǟ�����[s���N9�P�~��9,.L>GE��~Ͽ���0ј�Cz��T�?�eM�U�f�3@�π-�%8���4��%.qr:*ǉ�E��e����魟�D.���j�\���Ɣȴ� �t�u�Yd���K�����>��Q6���+��t���->;�$K�;�L�����K�F����9�km�Ь�PrI�F.;�T�� vY���Zp���c�	�O�MP�1Fu��i�v��������M���$��8�~x�@E��V�$�)�";�j,'�@3��}C���,E����Y:�Yg������S���x>:+�k0������Rc�gw���g2j%��#&j�Tn6OQi�j�e@�)�k56F̂�L������L�D��ꨤ1`Ek�J�)���s��ٱ����Ό�������L�J*4^�ϫf�b��m�k�#��Se�$Ш��{�?7!��
��5T�z�}��`�3r�O����n���՗��S��Cr��<0�tma� M��>؆{}m)�66Z��z�f���	Z{�.��V���h���:C��W�M�9�Z�Lb��K��FgZ=I��*Pp`��jl���aSU0�*ʂ��Q�Zk�����f0fx#&�������:��aC��M�]3ZX���+oQ)�z5dY�T������v�b��n�[�۶u`۶61UJ�sj ��D�T*BZ��ƀ|)�=ds�*T� ��
�^W�b�t�t�ij�AN7x����Ch�O��1���hm��#��u�p�7
��I��A�H�eޠiF׎*��׃t���$�kp�~�)>^�뷴cG� rE��p�~aJI����N]'Oj<�TtyN���zk�W���I�D2R�K���S}��	��x�G��"6���;���[d�o������
��)�TbH�#�ᒯ��}&�1�Z�L��:�P���r�zi6t�Q�&����D�r@���\3p��<F�m�?����Q��6�F���_���ہN��9ex��oWS9TK�/䳢1��C�:q�3p�%'HD�kL�z���]�ឿ?���>D��i.��-"5���1>Ǝ�a�~��7�]���PPo�[���'wa�'H�c�����z��M�!(�j�#�B����g�V����i|�����5{���J�զ���)��$�Td���L��$�� S�uIW�R��C]�NL��Rcʉ)�iI�)�T����\���>/�7��Ĵ��C�i>��K�x��F��R#�|UO��r���i�ͣ��S���+2-��\��JLݎ�XC��_�a��a���1���:+�T]y�+0M1Ǵ�;�<��(�#3�	�4�z������Q<��)0q�Qx���`܈���mW�����=�>��@�n��2�<�Hs�mìg�bӺ�{
��{n��7q��1����=�.�CO��t1�Smp։��Fk=�/:-��ߞ�	�v<�����!�Ԅ�#ġ��'����q=�G�kF�d����5��C}H�u�ķ�>W}�D$=�S�Ao� �y�}�utJ����q�A���>D#!D"a��a��x<H3[(S�S*!�b����T�>f�Pi���r�|��๷���X�HD� ੹���q�� Ǹ�\
!�S�y�O�iH4�
��l݉�k֩f�La�+K�e�e�����k6`���d1���ĹT���ݗ��������q�a�Q�eR�׷?��1,���7�p4a�)�ш�E8��F`ڏ�'4��뾉)c�*n��|V�\�ǟ|�d#Ǝ�1cZ1vL+2�,"��a�g۱}[�87�7"a(�Ǧ]��X�h)�;ې�?�����^�pHA=_�T����.f����4�
�&�b(���)S�;��N��_�|H�m���TY��,��#(&,	��T��R�02_��g�����1�"tww"*ᜳN�-7]�暸:���O/��7V��o����pD��j��S{��:����=ܔ~�k��j%F����͗-uB'��2|��W�l?��.B��ZG��Q^�!�,( �5��� �;�י� �K� Sj�hlH��3[�%�A�P��3�����)�7]B1�n���zDk�;���.�R�|
١��x���u1t딃��n���+��C�$��&�����#���4ŧ�cy����V�-�FZ�W�P;I�P��ʔ�&%�lei�zQw�G$c��g�C��Je�(��(�,�,aa&JBOss8�,<�¸&{Q�����5��f1���hO+fCV�n譆6��1���B�~��6��M��3�F�a5�Q�Y�qB��z�����D�즱"����[�H�4Uh�fpVs?4�6��z{V�N��6lK�?����P�LJvI"&<�r��1���+/�
N?�@�GT�&�)CS�kp�����u��Y�n��2��?�4�
N8�'���d)�W����9�-���v��)��>H��ܽ�ֿ�U��
L�v0�QM�� ���b�����Y�:���y)�2��j̨���<��6'8��7F�C]�/�T����)���
*�s\�	���&��
ZI>��G�}j*!��!�/HS��v�r���P��S��>dHgr��-�D�]�O��?%	>�\�rz�Qd(,�s^fB��L���x4��d���n�F��B��HV��L��sPFj"���5�Wb6���:��ak/[�OVnB�`�D���!w8_ ��@�U�?�Z��C�iM8���iL�vR+S(��Vt�<3���`w}{�����g� )y�%M֜�V{h�1��zoI��#�b~� �B�q�Q����0��m���>e�3���{}�Lz�~�!F>�!���'٥,Lc̾g��� M����Ϭ4��L]�kW�mnj�I�PFSo~�N�k�zш�6b�C�pa2 ��w�������$A�֎̜��z����/ kD����7��b���R����V:����_��#�G�;��C�?z=�:��������Ņ%���@��H�`H�+a�p�PJt�#C�7dU�aj'�ʴ�<_q�6��N��.�!oY�i0��$~���Ѽ�nu��LL#���ȧr����4B�ω%��lZ��!���}hN&ubڡ�\�rD��bNLy5�]ek�E��H�h����е�;1��� LI���4���
T���H�U^ ��(��(��#��K��&ʥ��Ĕ:�{}�^|eX&���%�s�!L91��ݏ��'����B���}�u�
��Q������� i��3���=b�l}?5|�}]�r��5�7^�-~�h��z������g�F���EFi���x1e�f|��Gc�=Ǡ��>��Y���/���mEa��I4�hA��H��t�e3+�0��T�����	TȦQH
ݠ4���w$���$q�䅯njL"���QJ�nL�p�TY۠�qe6mK�u���Rcz�o����fěG"���`j�������N�Ҁ��������[#�Nw� ��z���W��|�NA<�z���?(�L6/�xo�{-9b3v�p��$4�G����m�����rb�����D��C�Cڝ+��-1|��O�ۮ�F%dz.m���'��׿��{S��477c��m���������%˱c{��@�PD>�@:���~�2)DC�1i~���q�ɇ��Dy�<^�1���w0�%p���w��&	
y��t"5؉�Ӈ3O:w��k�����o���zc�b̂M��a̸q=�U:�#��H�;�\7mǆM��j�v�Z�=���ˈGʸ��3q�՗��N��˸�o�~��\����p^NK%�MWHR����<�Ҭ�\�*0�n"5���������`��zV�*k�π�XB����D�Չiޫ�Z`*����n�,���B�u2�"�5��4T�D)�ո�R�4L��!=�Tb_A�RX�
0��N��Q��4D-�1GsN��&����2b�O���W�>��a)�Y�YGT��}���Q�.�-�

�L1 J5��%�W�U�I����l��p%�\�>�_%Fc�bv$T�83`bEݍ.��A�����h3�h�5c��}�S0F���oP͎ܶ��E��* ��i�T�߷^�uH���2VV�~�kxHS1Ap�֑_0���ʚ6e����N���9Q[����1=�z-՞V�)��D��Kr�ظ��:[$p[�3�sWt�Z�jG��Y���aw��-��g�o�}Z��_c<# ���^����>�&��D��/��/F(��8�G�<:Ŕ3KЁ�.�*ݚ��N��4��Z,��r%���\�N���%���SP!��`�xY�P��R}*�E���� �U���������) �+��!�i��a߽&�Du���h��4U��	3+�Ź�eTdT�^������ȧ���{��ܗ�d%��{�Y3lsa��R�Z�$��t��!?�\f�+��6��R���,�2C�� ��Mso���=T��z���ޞŪ�[�n�v,_��?ۉ��+gz�4]zx(
�L�b5n�&�j�e�}%iHUW�6�-�6)��ԬN&�~w�Y�}����|��W�e/�^A�0�~��K��,͞b��ܨ ��AL��'�sN��|>e]��� Sx�w���Kѝ���'#��!DCQm�Ȥ+����Su����ժ4�̙b�R�+0����gO�&�JS��&�ڬ2�[��e�LӒ��x	N�b�LL/8����o@.����d�@�����r ��O�����W�'�o��݆��Y��� �Ӝ���    IDAT��#�w�_�M�ۑ���!V�@t��i� 6w�Q����3ݠځ�DU/��i3�*��Ma�:泫�ݳ��{D H��Py%r����z�>A7{���.�z���V~S���`J,�Zk�1�
L�1� SjL����R�����v��v�hW`���ĕ��Z���#�6�J����%�vU*oP�o�� U��_zi�&>v�����<��e:w�>�����hmi���3O�!�������~�yp���s���-?P'6SBho��}Uv�]_S7o� )U�ڻ�f7DW�f��<���dӈKLo��"z`k�p������F��G��|H���ڄ��u��{pO��Z|�z;u���PE@AJE@TPT,Xb�����x}R�)WMrs��$�4Q	(�� D�����af�̜���>k����f�G��9�w����k��מ���$���ݏa�
��Y��3�\�M���A)���ʒ�����j��2��wmqƭx�K�Ļ�r!ֱ yBv��}3� ?��d��V	�?��f���w����{�B����M(��Jj�̥D�Vm�P\0�[?Ƈ��m8��'�#�X�f�����W�'��Z����`G�8�iA���O�c��Qs�C���v�c��(�G����pI�\[F�t�z�1[��z�m�kL@�ڽ+M�����g����Tū�+��k�Q�;�c7g5�ʹ��@��i>'Z�l�0��X�c�ن������L?���p�w�?�V�|jv�Ɣ��+K{�\مq/.:�$�ݟ�3%Kx$e� ���-��k�`������Z�~�u�a���b��#�e�&m|V������kw�-r���0t0;S��n�矍�O;A��|M �����߹��z�ˤU�_j��
oaJ0���7��͵���;��^�`$qn�P����[�5.��Y ��zLC�K`*�9��k�^��J�t�2�Aˀ){5*��c:��\y�?���0'�1%0w��.�	���Lf�cj�5�>%���?<�������zU�&p�)���WF�����ul~�� �1�֌/K��ϒK4\��q�K��Y��$8���ץ�q#
<ְ_�Ś%�Dn�J9u��Wꉌ��p5� i�;IgԡXp��㶱���9-8��COcx��,��#�?0M+����z���'��8'� �*���	S1�l{�J�elb̩ѣ�&@̫��)�L���&I�0�����L�ɏO���ڋ������챵��>�
:�=��1�,#7X�L���s
���q�)�t{v�j
�w=��G?}-��C蠁��f��`��Ӟ�=�0	�q�*�q�<lמC�ٞ:t;��L���8`H�_Z9�$'�Ɵ[H}��.����̈��{�/A�L9hq6�M͍��߄�q�gk�~��8`�}��xƉ���M&F�WR��i�n+L)�+M잢д/d��љ� Q�r�v��+Y�JĆQ���6���㕯����t�x�M�j��`+cM'��/+�7�(�;�A̟�y�Q������/�};�11ɳo��lM����t4��~��JZvv�������p�g'{ڤ�qu�O��y�>�2t �t�g��zx�N�g���Ӵ�d�L�?Ɨ^��nk�QG���>�H��%��'��|����)�c.a ��F��+���~� v��0g}���?�g� 5}<|�����dl䬘�-	")s�p8��h7��'g猩!͌/z�ͅ��M�S9�ӧ�XD��� ��h^��S�o=�Ȓy\R�]���b5%|�:=
3|�$x��)��y0`̬�qܗdf����l7>}ōx|OO�q�(VqZ�{$��XF^�}*8��2L	�C�J:w�[P��<;#��E�>�u0��1%c�9�k�1hq�Z_�̏��cҨ�W�+�1�L�g�P)�afe2�;w��gQR^�f~�n�JY�$,):㦀i3t����w�nIye�T,
�jL�yt'�s2�����T%�İXL"��9V�̕��tj��K�9����c�x S�{�)`�Ê��+�|�JC���/</z��rhe���|�
|�_��P�H=<���?�G8�Ѝ�3K$I��ʾ�T$��#��0����w%e�捷����Jr�+��c[�?|�o�Y'�˅י �ɛp�7`0iȕ�\�T���=%����?J	vނf��&7}���'�1q+�Q�T�3��*<����� K2Ș�u�q��h-�k؋�9�}�+q ��e�A~��e�{R��g�>B0PH��a7�K�1Iy��;��E|��{P�ي��zE�G�q�k�\�A`�!����� �<�n��&��מ � ���İ�*܊�n�~�e�a���O��K��/��0WG�6�範ݿ�X�!��5��}LzK8y���;_����+qa��Q��i�d��� �8	�]%KS�����!%��|Cnt2�Ӷ��^�ͻ����	�fgP�T0��w�N�<-��;Y��faѦ��JI�]б�ӕs�]�VK�
�X5�+����~_�Q�I]?�ba��f��h4(ɳcZ���2>��W��7܍qi=�eV%��HPj�F�%��g��Ǔ>>�H�%�%0����*�9�h���a��OP%���ۻ����:ed[7"ߨi`4��Փ��7�L&���j�����t� _U��Ӑ��� SJNU��Ę�:�g9:��13��8(���T�=~Oj�Y��S�Q�c�>�.��k�oN�X���`���O��59 �ڴb}��cP����	��x'}���F}����h�̀�&t����c ��Hn�����ōAyRט�<�>�J� ���gDfXO>��!@g%Y�\I�����8�_���k�\�q+�"L�M�9�K=i�� -���@kG��,{��|k܄ӧ���IN�8ˬ�gMu�����,��u���&Iw:�"�{�%TS2�ueY����'���*��&��&N;�`��u/�1�fPgAм�-y�o�����	>q�5���D{BÑJ5��Xa�b�:ս9T�r�,v�p%��l�G/4-��u�L):Y(�y�2i;xB��V̐���Υ4s&�nk�	M����Ѡc2�J�@��d���+�k����k�أŉ���N8[�O�^U]G�?�?� ����s�7e���y�:P�W�w�a�J�=�$ovu�2�K�j���{d=��9��(�Eʬ�� �	"���
��#;p�mw��_݋G�܍�+-�3k�j[�4��tĎ�̨T���
vl�`��X��o�B��s~��E��,�g��8�M-�/LU*�F��We_��ɍɂ��B1�$5�b�O<�v������qg��*�;�8��-/�a[�?hk&^)�8�y��O}�z�rǃX������RCP4�JR����FpIG㣟l�W�eM�������[Ʉ�3Kg�������pB-"�rľ��f�����Z[�RnB���x�������R����&�YضH�W��&-��A1�+5��(	b��v��w�A��!��n����߽ �䈓�+<��w vHZ���9��L�C��������P
%��P!�27�!�e"{�3�n�8,�c:K���:c:`��`��T��zE���|����쓱&�p�ie,�\@s�"z2?*�ȿ��>�R��D�&E��2���H{�\@g�#W�\�S��K��2T�;)P�A��T]ci�����\ys�(�˭�g�w����ͧf�O	U�&W�1��g�������1��3q�9'�T�2����ӗ_�6e˓1�������7����8W��b$��1 ��������vƏՄGv��Wހ�\�C,,q�xU�[)M0�/�m��G��F�����>��~��?ވ��w0���ݍc;X]ZY]�<=�>�1j�)�Ju��yt�Զs�%�]i��](�$9^I,[)_ҽt0��׷&_�tVQ7��|�{��xΙO�:��r.����C����~F�^F��[˯�_j�������ן��?{���#_��� Θ�ަf��f���\�O���;�Ϩ17���sTZ�MX�����n�x�Q�@�w���]���zL���R]�喑�j�訯J����+8�x���n�K֟�J�k��cB.���Q1W�&�5�@t9P�g1�l�=Ms���Bob�tfn�{������^ۍV�N�߼�2-b�X�?���a�ID�T��\�������xa������?�����?�\e��������IB�J=�
�;r�|9�Z��2��l+��+cX*	���L���-Nr*ΐ��/����q/Cɴ��n�qҠȊ�P=�Q���J�_�6p`�[�<�\yɘg�T�	c,�����ʬ(t�.�:0�Y���H�(7���c�p~o��y'��]J�Xܐ�^���
,���F�˩�8�"ɯʔ�F���%my&�J��I���<up��ḱ)��@�w�)-�,��p�L��l�|їEIv*F��jk`knh�H������ՙbOtzϦ�%�7�g��q)���e�)@�"�B�A�@Hy0:@�~SIм*&�7����CksS�_-@S�Aq�fFitL+�Y�ݧS+��I�r�O�f�����0�K�k����	�}�:��e/�9���b���%�y�_�����ū����1.NdN�e�� �do,)P�kiV�h�5�^�,�X��y��otm�h*>���&,�KөB�>��P�'u4��kLo翝:��Pv�c������#�D��h�ob�1��*y�5*�~�!8��C���C�i���4g��^��'CFAZ��3x(�i�W�z����dA?� �L�Bq�
�eT��W�Y��ɧ���[�5z���p�3[۔R�a��
�xr=�ݹ�kh��hu�$Q J���Þ�bZ���U� �V�R��7�����M"��L�֚<�R��S+���J�������3��N��p�>�S=aq@̂G�]�w�� 2}z �������6��\�,�7g`��]�
�&n����b��������ϢW�J^�sZR���W�wd��Z�h�wꈔU��[8�")��SX����<L[��~y[�<��]�'�Hl5��RʵP���%<�~óŒ05�Af�V�>�{L�c���.f���lU�J�z^ZN�Luo��O|߾�^��j�+U�|����I/��L��]�r#K�sB�96Iy���Sp�阹[���z��J`8U*h\Ke8��N�����������*�+���\y�5� ZZٵ���E���N/�N+_��f|�@D�<��#�V+bL)��+o{������zL	L��C)�S{��a�\QC�M�ȳ���'�>���$�3�%\v���ל�������h|�3_×��]�j�8h����p��ǣF`JF��Ƨ?�5�;vp�����-3x�k.ƅ�93I���gDe+iʶ�[� �2*�\^t����Wތ/|�;XX&���*l��0���������&�z�\*�1�>�-|�ʛ%L�+��!X�ceu9q���K���h�g0�����#�_B�Lf��uWN��	���G�P��E=sE�Λ�9���rn��T�/����#��-�h4ؿX҆eғ/�!��YL��nĪnI�����S���$��d�:�1zr��t;���Amj#��b3��%�Q=�3�(�9�q	#��]oĩ��h�s�84�~���� ��W�� L�SF8����hȱF�Ȑ���p�}����sɂ�F^��1��6帘5��\��k�㶪��&Z��2Y�����\&I��M�ݩ���R<�G,4��~�F\�������̠L��	��Fsy'��%������e��@Ȯ�߷g.q���*nz+�L���s%�a1��ve����n��(ַ��_$3e1rL$b��@8BFG#���EUQ,Y��J��B!p�҈�?�pi���A�����)�����0�1�!0m��g�調�(�Y7��L�JQr�r�,�F���%0���QJLØ��`�"�1y�5l��Z�j��]|��G�e���s����Mv��I�o\�l����eP9��c�т�L���ZiFfU�xW =F{4Pu�X�J�3.�u8ɝ�>���ä��$�>���4�cԦ������J}VH�(_���G�U4l�(����INDz�pE1)3���5�8�Of $�5��Jd�YYiĄ�*��\��X�Z��K}Ċ{?pX��&��T�儚�NN�j�R�2_�n�x	��G��dݖ/[�hr}jN�y�c{k��c���;��r�u���u	!Y%�����������/߄��+��<S�wʳ��$�^�X����7��z;u߶����^����߄K!S`I��I��:g���� ����nv�M��_���zӔ`43���$�>2�x��G��v0ls�E�d`�~~��nݤ�m^7��7���#��M5}M�'{v�	.H�����5q-�����9��!�ή����xV(6��gD)�^��1�֦k�zC��A�޳��KkXkv�1�6��\R�[��<��+b�<g���b>U;e����ٙ�����%Cʘ	9�%�8���i�Ek͙�}��3�P,�9�a�ggqβjk	E��D��I�g�9i�c�6f����e��}^u��8��#��M�F�z�h
O\�p�-���Wބ��ߍΨ�!{5׺j��R�<+tjz�7��P�1���5�i���g	����� U�F��Lwe�PD�8��,B�-��B�&�ʅ.(�=뤃��})67 <a�E�ؠ�}�F���������j�Yٵ���͑��/Rz+n����1 ������#�r)�l�7�yL���{0�7飗��3A�L3�.Z�\�M��<�ʰF�2�U����z c�P��F�R�z}*�\-d* S��L2.]]؃��%t�=����Q��ŤZ��� ia��x�R�l�&?�兽���t"`ʂ6}=��TR^�n�&�́���h������c��Y,��N�;^s^L�}���1���G?s5� 0����6㲋��g�
+i�O_�'/��AE��ٙ���|́x�_��o��\&c�"�[0Ȭ�
�ra�����k���v������P.�Q-��o�0}�{ߌSO�*)o ӿ�����Wnĸ0���X��+�:�"?�c�l��|�>bff7྇��܉�w,k�L��p�a[p��XXX���{O�YS�4�QD�\E��L�`&S����Zk(�X}e�r�]]`�	kA'�2LLsE�m��m����&q��e<�㘐J����Fٌ(�)�ѝ���ml�D`�>є�,J�x�룛fs�1�8�H���C���i��@`�;^7�,�{g+t�s6�@�u53LJ-�d'��̒��Xm������I\��۰��X��An>
�Iv6R�Ѧ�[U4�o~	^|���pyU�����~T�LЗ�l����$����Y}{�I��>q~r�N���J ��6)b��+X[ځqw^��g�/�{�z�U�J��'�����}��Le1���$IK�S�x�9�'����q�=K@e��G��&
�Έ����(�P&��Y%e)��sh'>�$��7V�A��ƉLP����SJ�S��%��v��d���&�?��Ȫ�Z,���f��X��Y������� ������T�o()1g����'(Md��J�����}��۬�I_A�"�2�eG	0Ub�L�$��B�3�=���?&�%�>��D��5�	�«���stWu���V5�w���y���}F�x?�W��(ϒ����}	�b��c�FƜ�`̝��uG�����#I�k�L�V�Aw�4��g`τ_o���5���HJe�"�*KТ_6�÷ook$�㔰
O{*��͋B^�MR�������r������k%���"���+�$H�+��;�RAf(c�Io��.������p�G`�c?�@&E>�wJ����XƧ���{��    IDAT��G��Q�ΡP���8�N��Ö��1��w�X�MD�WJ�c�X����TW3��p���׊L��3�E����t6�NXro��`t��=�SA]��&��y�L���(S�ϣ~�a������lr��8`�ͨV�r��W�+]\�����y�5ʢ�J�|�w'ߒ�����E��m:X��č!��N����e<���ꞇp�CO��ؽ�D�ĕU�"�4p�#�BI�F���j���x3A,�ˠ�^����˩IxyG!S���TEA�qN�KzB[8���f��s��HT�Fj�l�>/s2���^��i�B���e��u��W�,�ԧ�|��#g�'����Z�|��Mk�v�^|�S_ů^�������s�hw���IM�{�b����@�4��+Ƀ�>�=�� ��Q���D[ 8b���Ĺ�͡t~.���TD�ӑ�F�<Dk�!{�<���p�	`=G���Y�꾿�� ���͍�������dG����ݎx/���4�+�(E1�jE��/$�3^�~�����Z����UD����'S�BƔ3�	L9GU�UAJp��ϼ�1���ӵ�SJyK�S�q�k��0�Y�� �4����)��C�.�c�muE��g1,���Hy�_cK`:W���ii�tVۖӑ�k�DLJg��Y����15P���4;���9J�~�I��*��W����y�yhp�}�P��w))�� ��g�����X��܊�\|�w��L�������q7�C����������p)�<d��x_�^�JٙJ���`lS�L�����o�׾}+v��0.T5��R��^�Á�Z��=�~�,��?ނg>m�d3����ȵ���<ʵY�#��(�ض�~����)�mÆu֌��_ ��5���O`0��c7�o�'[C���g��+�� @��g���s�"ʥ*J��d�� ��雑���)XI[͊,u����s���t1���@6���(h<قA�Vt��v��j	0A�|N�}Rb$����̊���j�Z�������*�Q�����vQ�]���*˨m{(�F���� ��^R"�>\n���u�m���oG	��Y�e��T�8�I����yw�t��vG��J�c2I%�t5����D���&=:�8��y��p��a�%�Y�{���R<p$=4^/��b"����-,�,$�˴�|���t/���O�co���tɘ�1c��Z^��)��}�~6�YR̃���d�)�A���ϕ�}S�L򑑃+1��<�[~����I�&ņ�X3J��Ő��M?��!4j��)��Q��W� c*ջ�lA�<��������,����l�t����[$��S�S�.l;�-S�K��V}��vd�N`Z���:���X@:�
��O�$c��/-��#0�,�yC���Y�NA����\Jg�2��a>Wfa��h5)�*)��^G�Av�Y�h0~�L��D�A��Sa�dRs���9�2a�~g��U�G9�l慒R��pdɜ )
�4�1�<�h�I�(�֤�']���L�<ɋ�7�t[>=\��Cn��w^�K����H �^�w%��w6L��zq��mO#B8�f.=Ů���ݕk?�i�v�l�k0���P鑭w���Oj/�����M���!���X���\�=�h��)�!��`�'G)�&(&��Š�������K�;���7��Ĕ��8���|���+�ފ��4J��R3��t�2�!KT3|��3�7a3Ղ?�S+��^�}���>���w�,ܷ`�GK�����g�E�Hm�^��3�dM�s���X�I�f�(��~�Mv�跛&[�1O�]�o�&�+s��Jؼy��f���[6���bf�,/�8x���xW�>&GOi����s��^}�`�R�<�S���V�ʥ���..c��e����o�� ����n��Ǹ&�j¤��wUE1�|m�s��pi����#��H��(��������-;����rj��M�T!�7%���[�K�1�8�^8YV�{��Q��}���e(	�ș��lI�C�?��XW�sO«_r?�,�P��jp3/��{����>(��G��ѝ4ПT�+�)֊�G���;���}
����@��m2��|q뾳.���3��e�J'q,�Ә�f  �"e|D`J�	[��&=t[;0�-b�\��'����ٜ<{=�������|��@J��r=)F�}ƹj�����^��	pLS�;�Z{�'w���_<�'�t��ծ��R��O$���E��L{�����.�6���c�e$��y����̴�%þ��X�ə�9�
9Ls4�x��Ԥ���@)o��'Әb�2&d�l丘�����s��)�I���(��`�R^2��b��N�L��uJy	L)Sg�/ӈT�)�G>�� ��M�t��HnI����Ұ���2^{����W�+`���ݘ���)ӿ��U2?�80}-����Qs��G>�-�ɘ�P3�3�r�_s�y<�Y'�����������̊gV�G��}<
)g�u�N\��[�ß=�f��5&���閚�R=�zdogw	�����x�	ĘF�/>�5|���a�#[:-֍}�[6��W]�K�?U)��K]��ǿ��X@.7���n����:���,`��?�����{^B�<�)+��V���F_�"C�\b���H��=4J���x�Gw��`�?�P��Р�V��1�D\�6�tm4��$Yg3Z�אe��8K�s)k�iIkT��&��ob��0Y�9�e����-�~ԑ����'3髇��3j��0�sv�j%���U�}�� Ӭ�"��%���צ����U��UT�HK��
fõ�{恠������1雼���Zq�C�[�Cڂ����\*h~�
<d�6GV�-g0%����Q�P��eA�����
~u�.,�iTG}j�*C��}��^{����}\��3q���0;]�T�k�?9�40>����MNk2�1'��Y�� g�Ȫ��c�=��k���w�'w>�g1P��:=W�x'���nv0@�o�K��I�"�LT�������q��4󣱜��c�w	��5�T��j�����)=�P�!G_�!�MJyW�[k*X�5Iy�#w����+�>WSf2������S꩑=�`�� �d��>$�	M�~T���N�ٱ���M+�!�WR�����j�$�~��z�n�i&����2f��C
3:bOi�\B�^���5�&���q�h���d?�8+�#a�;��b�������X)#�g/MW ���SS��$��{��^K$U��r�c]�%}��e	���W�٩�R�SK��Z�e�_R���,�Yh������^[�*F����]I�H��4�l�k@cr�+���qI�W�����0��4�;�#���0��n��x���-��n��rC�Ҍ�ȌE�)�����	|�+7���0Ԙ��z����X/$�={�z��'��kĝGc�'�"���/6�v�ۦA�憧�_@�߹)82N����7z/���hf/����ml����h���S�$�-U;��t��������3�d�G�T0sA�"`q�n7E#�`��5���6m��y�sk���T�.�E1P�Qj�2���c�L�8�n8��3Jz���<�s��blD�FW��V�A��b��j����;T��Mj����.�*x'fm���[���{q�ݤ��/����=�.��go���[6a6a�$�E�e))�X����~�{;�������A�(ފD`�<�q�o�G�pƨ�c�mī.~6^p���L�0a����k;��~�V|�;?Ǝ�	&�yt�%�E�r�g�r���ª;����c���nx�y�͐��X-��LbJ��s��>M�?���,�d�N���;��*����\|��$ϹQOϑ�c��	���e��
*f��*O1)�\I��Hd(Y�f�&���i�X]����XuI+���߀���́��C�IdR<
1~��1�po�,��2`�y�r�8�V+o'���l&�����C����4
s3;0LF:[+&�2�^9E�1��`���|!.��Ϣ�a�Ӽ���ɔ��zL˘��U�7ƴ�!�<�C4�bLi2��st��B4����8�l�1�>�Ea����
^�Ix�+��)MrO���GnO�IƔ���&��Ԁ�Q���~�����>wƃ)�>������0�Q���'l߆g>��}���hܩ���8�R�����~z�}�ƍ?�C�/�/ӛ�L|�d�t��N�>�d�8z�:���^�SNX�R��u�����W�����I�1��ǘj�������p�AE�\��=�sW?�O|�����5s���]���'�i�-�����O� _��{ȗf1������ц��j���Pg	(�e.D���a�s�8�
(r���ʥ2����f�m��n���̥L;��l�	={����I%nB�|hO��nl�,�I�.z����ݕ������*֖�Z݋q�%���G�N ��,�Qհ��Ґcs�֏C��Y�[�@��<�DO�Caj�j�b�+�6��}�4�P��a���Q�tI� \ܧd��Q:��lI&��!eϴ0��ϗ	+�r�i���v0aE�%�%V��<l�7�e��Qk?d�U�|YÚ9��\��ԉ3P9М��C����M��(qL����z$���d�L�ɛ���W�,j�*����4<���.�������D��������Z�M7�`��*C)���^��������	8�fi�:�4)��&����	�5�TY���"�W�����%�lo���*�˫	0��o+r�?�
`�3����22v�a!0]ZF��Ҿ+�j��������0�)�h�1e�룷wY�K���4��'�.���v@�(��0ß���5iɮ�Y���y����4�����H;�u�$��CY"	��u�*U~͌.}�8s���+*�55�3��z3�b�	��^���ݷ{�{bJ��G{.�T�b���w�U��%��X��	j̥���� ȓ˞y /=�d��Y���g�L�k��3��6��پ�i'�%;�R�8�&7�֒XsK+���fIF�� � ��d�7O��jZб�#(�I�^���eGϼ,*�T�/��ȹ	:{��"��%\��S��K���G�k�`�9��i�����W�n��x�q}T1��2*d��9ػ�"�"�h,d=F��?(uo��Y��5��,��W���H�M�M!�3��bw�(K�*�?{VJ����b�������x�� ������l�v�sy�}kGTXŴxN����m��3w���8l�O̔����#��R:�s��l�����/5��/Bʅ�&>Vl5EG���2�m�	��g�W�0r���c��S��w�q᚜-��;#F5eƲ�q�8�Mz�Ӿʤ�O�T�����}t�ӭ8�a�=�\IF�1_ўjYG��Ĩ��F���xƑx�%���'l4����?;z}����g��p;v,sx�,Fy*Y8�l�Uv�${c�  i�BT�l���R�O� 'J7���g�Ť��)�_�c-d����$	�pY����	�!��>��U��'��H԰��[-kfH#22�T�<�b��R%��<�9c4��K��
)Ek}�Hͷ������gP�N�X�� ��wc©�!B|�s���Z�xz*r��Ġ#
5#�3������J�+W^�����_/�1[)�:���w�̏F.�-6�L�ʛ7W�d�9�<&�
��w2Fsa/V��-g]΅��ϡ�~�r%������?6�8c�j=���KyW�ڧyN(�2`JP�2���@a��j S���c�^Td61�[�^x
�z�L��������SW�+�ތ��:l;`+^����ӎ��]o�Ͽ~���ZLFS�K8���ј��js��w����eLz-���`�A�p�~q��1GV�TF����b;���ѝKxx�v-w�ۘ^'�BѬ���b1/n�k�;l/���7�=�s�q�:��ϣ9b�W�o��Q�F��&����E�;��[/��������� >�ٛp�wnG�=@�<���Kx�[_�=��\0�A_��N�����<�9�j�Qa A���y�k^��Q�َa�>Q�	<|��7�a�9�&��d��jL��<��Z�d��)��1*���M:;� O��6�1m 5��,����D&�a�jT������N���J~��2j��KY2
�8r�l�ݜc���b�N7�!J��X,V���1���z�L!_�������&%c��A=l!�َL��S�L�t�y�t�? ��L�m�*Z�0�)�Q�W�q5�Whl�-+L��D����[��Z���%;��K�h�J�JE@OE>ʍc,��&�	�7i�n��\E�m�u�!���k��Q�V�����X]]��Z�%TV������Q@�콣��F��q�R��Ą�-�.�y&,�=OZ��0~�>�-T4����J�9��e��*d�K�	R�b\��i�j)	��1X^Ck�R�1s�hl�().�)���g���k�|�)�V�l��˯)Qʛ�d�x�K~�dW\C�t��.� O%�*�d����]�N�l���>'�*Qsfv�����aK��^�O�W�a����ZZ"�՟QPS'�s�KGR�	���X�#�\̣B���s�u��kP�a�b}���@��L�1�74�#Jx�&��_�\"Uiv�H�v��5�P�Ĕ��W]�k0e�7��Jm�!ў�#w�¥}���!3���K�G�'Ya�#`b�&S%�>�Mʍ�
Y]�`3�D�͸'}�.�uH�ȺÜ)�x�&᳘`?�טqn�	+��,hJN��l��,����a{��^T�M�&��5�٧*��m]�	����H�������oފ��t�&��Li���@����B� ��u+�ؘ�nRS��|>)&���W��R6Y�b����_j�$"/����G�M���^��0�k�"��wΰ�kɺV�Ķ7����z�� k��|��O�1�ﶟ���FTY���U��E��\b]���ħ��\���hl�m2제��ˎ�Yk_�Lunv"�X�R��~wň�R��!�r�miK���4 ��������?8�d9��4Zv���=�G��jD?[Kv]a�fc/x�b���ę�|�6:+�8���矆W��98|?��3�G$��[�6�ՔF���U\����[~��^�IM����&p��.�Dz.�U|��Y�R$�̳;���J�v�R�a��W�w{NFlX���}��F/�d��<�ݥ#��'+�c�H�5,��������w�7#�z�Љ{׻Q!؍�d�f#�p�I��P�68�\��נׂڇ����B
�G$U�2�HFe��ֈ�����1�T�1������*��Qg>���V �9N��w�=�c3F�^G~�R޲S�	k�3��1��1����;]���H)Q[7/`;�RCcW>#�	T㸘r�5��;�ovu�0�+�r�"�yR�k���VL�5�� zL���uQQʻ��\t*����$��l<NNi2�4?�����W��u2?z��¹�[�)�����&�ç� W�`X@cv�*g,�1�s����%����h��Ԝ̒��)�b��p�D��F�P���rI;[ �	�&b��S�^�qoG���w��glU���!c�?��
\s�L]���1?��e��7��r�|dw�������+h�k(ьh��g�t��a�a�P(��9��=0ě���Gs�x�e�`�&x����o*j��^n�	m�(՘���3�*r�U��I��1	���d")���e�L�� ���$F%W	5�"G��Q�w��d�t�46O}�IJ�d�]L�M4���E���O��[�Q����ɆVZ=<���o��Op�?Bo�j}�q�	����q�A�Pb������>~v����wᇿ|��zL�e�%�>K�o�g�x��X�a��H�
�L>��� �����p6���ʤ��^�Isl[�ZpP�\DU2���3�    IDATU��#�\�E��VP�U����	��;�ɳ�0����N�9>w��n5�]��&95�� Ч�Vϋ4�h�^�f�奥%���*���qW>;TCc�H̫��u&��~+�������Q���s���hӳS!�O9�\�KR	��/��;)!W�C����Li/U���%�>&�|&���Ŵ�W��s��ڼ��0�q�̏Ș�l܌�i�֛̏�wP���s���KkG}�c�}`��*I/G	0e`
@�+!��S�I>�'�^%�nH�U W2RIfc��-��o{6��5�A2j{U7�?�Ө�ӈ��
-�B�(��]��!m�&��,J��	Y��A�"������>F��,`O��̑PI�GJhL��܋p�31�O5(뮶�w��@j��	?K<NLv\ea�W�kd����O�L�
��j&�K��Sz�����,L0�ڇ��$����&o�si}�/�`�#!ו�:���{�DR�"I�,&�h}l�[�jz��!���q{6L���9x�������wK� �&,�p���7���%|�K��;�r�����jo`�0A��/�
�����+T<w�g{�YV&�8I�D8cb� +\04��>>[+��|$�*�f�c��R�B}7�Sh�E�0Ak_�,\ś?'�l�y����-��9��k�$�16b@���9P�Z���n� ��&e'WX!ŀ�~w2���yƠJ]�2Q)>DӺ��͸͋1���EK�T�L�kp����j��@|�R񉯍�ȡ ��|3�Mp#ޅ֮��l��3/�����>2^\�|�MZ��1[�iGn��.� �<n�&(�gSI����߁�I�5č?�9���Ǹ��
��0!S� J�%?�������y�(�S�s�'��c� ���~HY� '"rĺHT�Ĝ��̙�3
J�H�m��]E�����:�_mP�X�t�����(��YWo��C��<'���e��W�g���:(�B�����\�,�*�t`��%�ZG�E�z��Dq9����}���gШ��H~�K2���˔�^(@�t40�6Ř�u��@~~�ZY�|��n*&���%`����X۵hR�rչ9����%��0T���̏&�)��1�"�S��ȱ�ufZm[������<��y,!>QaR�� ���%��Pl��/>o����;`��ӏ~�:|��@c~#���~�8����T����#��7�z%L�%�+U��ǀ�뛕��L�����ڔl
nF5���L�2O��}�=���yY�ˮ]f7���5y�<���ދ��8ԪglF0�2����1��ѧ6�0���	��s��K��ƺm�;؍˯���lc�~�`�!ȸ`��b�:�K_x�=j�z�ᮇ���wK�)��U��SbLYa�K��JR��ha�i��^H��>��!f�8��h�6d(����ŵ������Ҁ�ÿ��Ӥ<��B�='�өj��0!���Ω��B���h�����z-����_��-ض?TU����n�IH�����?�O~�:�ܽ��u���^�3NZ�y����2�Y�7޶���k5�q������qn��	�ٗI����jZe9f���8���Ț�9Rv/*P�[����7d�4~%����n��-s�>�j�snYuc�n�ʂ��N2+�@N��&�Ȓ�;�$�fj���D�������%SN���v��u���M��,�ʠ=��r
,��ؼ��c�oC�^F�RD�a���=kx��<�cU��z�l��@�0҈&2�F�}����'W�cy�A���*i� /��8�b���d�9G�zL���gL�?1ň���u�Y}��w�=�m}����LM�¾	���O S:#�[S�����k��G:P�#J��k��'`�*��l�+�������n�G��k8ۏI�?�J�Ƙ�0fI�l�?�9�cI�;�'��i��R�����+�&쇨Y��tޕ]�����6F�8�Y�!��J�� `��`�,Y`Z쮏��a��h�6<���X{.�K&�e\_��F�o��02��ӄ��Y�>>�[���e���:\2
�g����i ��R��G_���@
/^����x�J��4�Ai�(���'��W����|+)s��
V�O���u�������(4q�)G�E�=�8�P��)E��$�V,H�Kg�����v\�����b��,���mc������%�.Ƕ����ھ�=d���I�&�!�
(eV�qTN�%�e�� }xRJXەޯ���2�][ӶW3�{�_Yh�ك�Wkc�kv6�֑�h��π#}�3����\�yd�:���^�p{���'�������ZO�Aj<3[�����Fޞ��Fٗ��W�Y�E�P~ا
xNޒ��9��ad�bLRg+��M֚Q�	)���,��3�)����v
�=#/�������1�=�z$C0�0j�Э�8ﬧ�瞌m[�
�%*���=Dl�\�O����o|7�r��
��i��eX�	$��ęC�dߐ��4��Q-y��%=��u	B�@}��DN�$ ~�¢04��IF���x����;�����s �ٽ�@��S�Q�c�H�[,fO�`�YZQ��/���k����F���<-\���V�r3��8��؛I$
\/z�8�)184Ɣ�^F��N������1�ǔW�c��J%�VJ��GX۳핦M� 92Ր+/�A���0������g1�l���k7�K�'_D}�z�8�Z��3���.�vƔ��L�k�0�sL���
'0�0Ȼ����M��L��6���oL;��1}�KO�^|�ZD���)�)]y?��kLk�����x�K��瞶݀i����>����a�M�u�
2)l^f%�M=�}3�V���Ӣ����yH�y�T�;�yh�[ٓ�%�B�=3k�v�����y���U�^�Ⱦ�W�7��I�W�6��W>���������b���&%L5f0C�3c����M�P����x5����m��Wh���Q�������Lm�.�<:�&]����
��̣�җ<���z	��;�Z���;q�7���ڃɸ�\���F��jb��V��K�93̊�o2��D����3Ys���Tߏ��v�P����0�a�݃��;������sE���?�q��	���_��Gu0.}���ܶ"�P���s���?����V�%��ǚ��q*��,�_���r[�C�{�\B0���Y�)�hc2�ǔ�a��q��!�*s��'KO 8K���B��D���.��1���g��KY/�
��[�t�����4�`J0dF`SKi��dz��
X+q�J?'�_���L�	����J��S�1���XN��cR>\�t0l��	Gm�E���9�<���h�]��G���߸O�؃Z5��^r�>|Z�������Pҿ�|��'p�����~&Q����xa`%-�����1�Ř�7oB���sc�	��!��T1��ubH�t�����Y�\7��ܴ\yi�R^�����aZ&�-h�0����`���%kf(In�k�Ұ�mӌ�X�$'�B�}7`cgu�e�i�15��^� �����K;ju�Rz�^�	���@9�h�#a��&� p�Iӑ%��oLnh����n_�tRĢ6�ND��F�Q�;���{��KcRB>�R+_X�/�4i'Fw��x�� �ޣ�0�ztf���cWVPsbn����+�U����VO\	�s���$�� 9_�um�Y�&�n���J1�d�kr��H���8$ZA-~gM?|�9��)��T�~�7�B�&#c��9y,��C5jc��%G�C����{*^r��ز>��)2!��g..�w�z_��M����j�#���b��r��4J��+E�L�Mg�,��S')���P�m�*ęv�RKB��L@���IO���9��:-�������/ט� �!���B���f�`K#�3�'�:�榵zKx͉6	�u�̰�:w���Y{�[d��¹��R�o�'dL�t6y��u��v��I�m����*q�V��=�a����Ґ�n�2a4����yd�6V:�W�w�>�����"���9��2�>ߝ�@�T�-%0�P˷p�3������۬�Y�	���)c2Y�GvMp����u7܆{^@����SR�r%S���X�8�|*0O�m���P�9��'��눕�1.���\��u�U��`C:�U���,i�m�@T�Wo��1<���Sȵ����*�|�\̻�5#��3A(3�_�m�h�S�W�PQ�1��΅P%،M�6w�*O��u�[T����J[yv�5���b�� !{���<3��Ex>����ۋ��E�q��x�U�F���Cҿ�ʲ<]yk�#Q-,�ffq�RH��+dLw/�ߦ'L	52�s�	0�Z�,�bj<�\��9Jy�m1��qUNR.�B`\)cT$&�Ϸ��`���%���YDH`�Ey�ĺ����3��*���U�w���\k2�4)�����+����v�V����g�S������g/��g����$�b�8&��?%3EPR��H�ߨ���l2/�4�T%����ƻ�2�LV��KG4ז1vP.�5��C7�����S׾��1��?�W|�_ ��Z7��i���.9o~�1�B��cL�#�\�C�%5V���������'��wG�.�-V�E;P�\�Y�-e����6��LU�8�ԣ��o�PD%�B8�6������t=y�I�����/��s�l�VF��۷��[~���b%9'C����D��r %���yQ0����m�~�V��J���k/�[_}�f��s�,���;�N�T��$���ފ����9g����$�(1 �T#�Q�O�c��wݳ�By�:�<ʙ;��GY,$jqx�e�W�%���J)l��q�����8��#����Ӻ�1yr7n��A���]hv�+5�n��4n�����N4jt��UX\�bR�B�1oV߬R)�27-���E�����A���$%��Ŕ�Ad=q�[,dz��b9�Y ��*b�WWV1�s��@�BC�l�
Vy�.N:j#���p��%I�='I�+��?�ţ��D���g�v<6̥�T��SM�r�B��<�+��{�U��)u֌C�l�lr�S��]�����W�+3�hlބ�tCC�y 8>W�S<��&y����0�{P2��'-��S2��j�h2��4����R�	;���3�m�ŖEbA��y�:c	[���zN���0���)yp1f����&+N���Vh�VS�$��7R'�:�2��"�]>��|dn� ��)�w�z��i�H�x�LH�$C�!��LS��e�>V�Y���Xϧ�
H��:ښ'���4��<�H\!c���S���	5��z�� �}��7�gf�ٲ�]2.���� �׎[�*�jT��ܘS��ǱE
 �V�+�!	N�>[-�p&U�2qM&�F�0X2F��4c�@��"0l���G3/8��x�[^���BU#�l���L�0gν ��\w���+o�ct���4�RuJJ*P%�d<`��r�a�h��Ո'c͍�1H���]����<�����W�Q�	uV�33�~��>�(v�+>z��ɪ퉌�R@œg�S�\���:���������k�}�K����c�= �]�%�nJ�kYN��ܨJ�����k��{�~qk�3/���Gh��Ĵ(*h��n!����[�/���*��r*%I�B�B�'b��yɷF��M��4Q���S�N��
��&��1�[_ŋ�?�}�Y�2k�1�J���gGU{���}�����7�;���+Ϡ<=��x,�sG���4��1�	�g���3B+'}��&_k��;�}���E1�e�o�ɿ޻��xV	�m��s)~��L�M��}�����A��EAN�w|��k�K�*�<"���#Y�4�������:O�LK�B}�1�L6J���$����-���E��e爝9i�=hKM}�����H���N,�9��f~D!iH�1��˖�F�(�*F���F�@~֤���ȼ#[���V+�1?UGe<Ѹ��݋��V��Q^7+uO���-���c:_�`�Zs�t�H ��rQ�i�Be\^����Z�Ȣq`�i*�{G�d�ĘV'm��V�W���.<��k��;)�SW܈����غao}�xΩG�ǔ1|�I��6:]�E4Za��[���5&�\ȞY��i���99H�3�I˚lU���b )�ǘ��a��ih:{Ș�w��gpӭ�"7�c$��	��#�s�xǛ^�#����N1;I�5B����-{���>{3���`R`��#_*k��h~�2������܌�{<��ܓ�e�����$��~���{��߆�=/y�i�	%���_�?�E,u��J(Uk�q4���}���3S P���X�b����šLAsu��2�X���b���'��S���j���{0;;��ۏ�����x�h߼�.U�?��T�=;���}/��N?�l;h��e���������nG���4�u�9G��L���W�� 0� ]B���x�5�}�Gou/�>t#~�7/�'oE�H$%�܋�j>�p��~��o�O�����0U�`�>��mq�O�g�������r�cX��5��}���.a�CӍ�0�xI����uo�b
�z0�T$�!4M7�ѥX�:ߖ������,Wa3� � @�7�':�`�����:���yUw��|4��:��{�i4[CL5��6�#�&�<8i2��^���_���XVѧi���n]�5^�d�c����*ZK�cʞ����
�7�@i�YگF�d�	L9z�enɍ
��bLŜIy���gSF�r���4?��hP|r	Q$C����O�VEЙ�O枛J|�kT�Vϊ}TV��7�e�MC���剤\�@˙+�)ev�C�FP�GL0�@��m�mp&_�-���ᡢz0Ĩ�ќ�H��X6}Mb0�	������F�&ƚg�k5ӏ�~�wSgNK&R)V� !u������^B�/��K�#��b'+��?�3l����o�@)ѳu���b)������I��N�������$?u�S�ߐ����@�eȔ�0�(���=gUĕX�a��D��h��E�����n���p�����o|9�:�H�S��,�<H��ď��}��4��[���Z	�I(�\��Z��B���5���s��um��P���
~)85 d�V���剹��#l�[C^6Vo[��j��}��/��^8�j*���2�z�������� ���o����(k�eWK88O�dqq~��UpK�`:�&�!VL�]���k�%��hƧ�7�qޟ��h��)ѷL=�~6[�a,x@Ocģ�c&�N�\]*-V*���<og��i�+#D�Y��p,6��ͺMޗ?��M����oH'X1w]��dJ����X?S�i'�W\�l��3TN�ҫ�X~͊�JWz���ۋ�}�z���{��Q��@�2��ofE;�w��S%�'_c�@�h���ge�$ˑ�]��SP�]�s��E�s� �c8[-���7��t]�^��2�8B���� q�oT$8M!�r�p�W<�rM�wF+�Ic�D�,�R���؆!S��� �6���L䤕�@�Xp��Sj*�tm�����$�<We��G��V�1��Ο�'�Tu5��[Bi<�+oK�����(�ظ��%�I����+���r�C>����Z\�S�S	Li9��L~7,�Xpa\`�6W-90�+/�3?ʕJr�%c:�S	�Õ�ǜ�ڽ�����ۘ.�d5�ۨ�[�����矄*I�l&��te��h�E_����˿�������w��}�!�+�}Jr!P�^_���]'X����f�d���� lqHğ3��ă˥�:HX�%0����+~���5���9������矁�<�xl�=�g�t�y�0����v�l5�/�ӛ��Gw�{?�W}��^
�ywQ�(��%?�;Å��e��:�a�ۋ�{��x�EGa.y�Tc�E&�Ƙ�1�I>C��N0��a�bH��    IDAT�1��{�.���K�z�l����)=z1�6��\��E�ֿ�yK ���b��[M�Z{Q����o�o}�ɨ�������|����4�����x�.Ÿ � _��.�}����~���p�}`�o����\���c�l�B;�������p�Æ�3���t:�����F�T뭕L�����J�a*���^w1.>�(�rz��5��H��xx7���~�˯�.Z�1r�6��\����W>���Vhv׃����5��e9	��$�J�z)��В�w	�ڜI�Gc�R�P�����z� ]��033��Sʵ�e�Ee��*e��f���)`?"E
Zk8dS��o��[���YdGw/�I��y�\B����v�#p�k��Jz�	:�VZ�6;h�Gxh�*n��A���&[*�[�Aq����Ll�����@��c*)�>�6㮼���4�$��Th
P�3[k���q1m=3�՚�Ay~F���)�k������lA����e��0O&bL�y �������� ͔&3�����	�rj�_=!�N�C7	��i ��tK�����uW�'��H�g�w�W+��x��6wٕW�F9��3sMU��6C�]�[���o�DZ�gN�*�D��%���!C��XwU�DV�ERf���Lpv�A[�@�y��p�s� fE�*�/�=�15Y A`�X�0�T���9e Ձ��]�W�=us@�`��2%�8�QJu ���-	�'A���o��}t\��ء�%�#k&�R�
Uj�{���Wˑw�A��ݵۻq��sx�K��E矆�3iB.�3�!�+������{W~�Ǹ�'�c���so�JsĚ��*[ۏ��!(pC�x/6�ɆEϦ7�i���<�����,��~J�H�\��F�����O�4�p�G�Q��9��E�L-=��Q���X��@Z����uC�m  @��Ĝɪ׉$3֬�[�8�M�+���_׮�a����y,qh��;b$�v���'*����IL�l��`YXt�U�h����mۏ��l���3\N�zQ;�d����"�_;�\'G#0��wښ5�oӰ��Zi�V��\x^x�)8t��T�������(ݵ|����݉_?�G��|yy�gP�����`�b�Z5�0�mk�&��S�_S���3�4.�
ba���eLu�x�8�G�}d��Q8��+��oH%�p�{��\��r"��B���3�\6�>�W����nR�I����R)�+c_�yW㳱3UJ�_��l�<?��ߑ=Ȁ0�J�#��T@�Vm)����u}��Zi�u|���Z-�.�(SY�wH 	$@ ���������~o�~=�9���}��y��}_�u^�y��P��y�[ؐf���p�L�����}-ž�I�t�=�s����Pǡ�G�XU^6Ҽc��Ll����_�mczt����R@�ߛ4*/}�)t��5�uf�GU^2\'���|K򥴈����o[����b�>�Y���E�Tb>�L�0m�����	B`J��h�t���,9�:ҝ�M���l���6z��8��k��o���2��'.�N^�Rؑ`MZ�U��Q����8 ��쒋�$��Y�G��~��U>d�6��~�<��dR���q��4��q�e�Xs�rQ�]���E��Dy�3��GV�K%,_��|�G�p�C���{���$���!�@H��d�3�jzm׎��V��v��vu����������S�;�s:/lۅ�6����I{��v%�9��H=�)���D$���{�o_×�v5�A4�F&_���&�*��U'� �������(��/U��wQ-W�(�!��_\~!.����AI
�?�y�t��K�ǧ�����?�R��:���n�u7���ڋ�]��:=�d��eK���_�"N9a�j��ͪ��<�:(	iS*^>s%t̶$���3e
θ*�a���b���&޶f9>���0� Ms�r+�cJ�D
��ށo}���!]tG8��?�I�,�K�
���7o��[����'�oi����.] P�Be��L�FA�*�	I9��*�0�E`��R�Ѿ�4e�Y$� ������Q�V��4��8�A|�>�E%�|�=�u\����νx�y���#EL��MUv#0U��.��'�wd�UT�<�e'n��)�:�F/���y@�y��*��@\��̉����61��Դ��\���LC��},=Xm�mL(�>SAC�iE�i�����1�����b?B�SvL{�ZcS2�����A�.�Ϊ������9��٬�S�|����g���P�k���Sb�W�H	ߧ�D*Xsʫ�[�N�Y)m��L'����HE�%f֜S��'�]�@�l��љ���R��Q��T�jM��������D�1�Ж�~��Vgx|n�o��N�V��nl�Mr��HI2�œ��j�
N��M8�	q@!z�Ȑ����ʈO�>�hG�;a�4��+5Vc�$�֑P�R�
��u�@��4�.Me	@�Q���{Ⱥw����
-�f��<yb���1�)T��&H���VB`J�D�t%�$l�t�����MoN��i�]N�.<+�%ىj0�yǈwZ�l{��_��(���>LT�Hd��t�$���
z�@�]9/�Y�S
��g;J�	��=�g4�)�l��'�rvX��#O>�εSD�;��Y���V��O��Շr�y!"z��_ ���g(tt@���ϺN�E�n�l �b�o����B9Ѯ��q������WHŢ��;RzvM�L��,��~R`W��+�O��K��7ػ��,5�vJ1�U|e�Fܤp#J�Kt�h���E�U{(OOajb=�[5fkOc���<�x�s�I8���0���.2��>��1�Wެ㚟����y��te�wb���0!��:��@T|��!!tP�쳙4���#g�ȳ4�?sJ�/L$��/��쥎K���0~9�Eϊw��o�~i� �V2K�#L�y��3���$�Fٵ��V���i�$_csÞ�rm�}���w5}M��o��,\2�b���U�c&|h�����_�ɬ1�E����N���cKt��s��f�HL�LS���r�7Y�/pt�_fD��(!�6G�����]z�d�tl
�rH��D�ʺ��ف����PYm��e2��[�;���Z��2Id���jǔ�G��w �n5+����a)D��c��d��Dk�|��3��GK�Sr�h�-r�Ś�^����v�|#���T��S����-T��-�J�4,���y�F�rb���묂�w�����Ϗ�]�v��~� Z���G���^eG�t�xR���n���	�Mv�"|𒋰�c0g��-�k�Ij��b�Ρ}z;�~�%���(��稧#=�X}���a�:�2��Q��ʸ�G���WŐQ�H��k_��O��/��J����G.�C�^���N#�`�>�-%�����ln`;��[7��.�zh�t�TĢ� �l�#NIL��T�	��pC���*��Q��c��'?���(Pє��w�>��~�[��-�o	.����c��S���a\}��ػ{��r��}�����A�g���&�����M�bێ	 QR.��=��J��.#�Pe���S,䳈�
-:hէ�x �����8���D�]�������l.�<��(���7��7�`q_v��xﻏB��z�v2S5|����=�l�X"�t&�E�$AP�@�Вl�8�?�N�MLE(�B��=/;�(ͬ��5=|��J� ��S��mD 1������ݯ\����#�q�>���a뫻1g�",^� G�9k֬���0�����K��`<�Ĉ�H�`�������շ㕡fzE��Y ��b��j�M���
0�������t:ȕJ(.X(�\�tB��8���G����g[�����҈���"Rs��+�ù&�2�n#1-b��//�j͑	�2�MR�"'�Oj!%Tb�	�h��_V���A�%�L:��$��DZhD�C�k(�5L4�aF;�L�0SId
9$���b,P���҄D�@f�X(M�_[=��%mS��3�P�:����U� yW�����pP����5iՓ ,��������� �jy��;�<1��>O��vn�>K�i��Z��bN���S�s'��[)vq��e���Z#�d\l�@h��)��`�:��(���~n�\�_��5���G�����PT8ȭ9\]=؝��,a�=z��+�B������hC��z[�h�SA�>��X���K/>��t�u�J�� ����z���4��n�~r3��4:���~$�E�O7ő�'X?_8�n��π����B^0f�kj7�mJ�ӎ�f$Q�MZuOYo�:��Wڊ#�P�N]q���z�i#	�S)�X���ÂWE
���l�� A����+ж�g9��g"g"(����}�qt\�s4}.^v��(�@Ɂ�����tdJ����W�`�\)� Bi�xi�Ua3�q���K�IZdy��T���Q�B6��N;�(\|�;���A�T܈EZ����4�Gb���x��-���y�0���]��D{��r,�C�
Z�`y� e���ZO�|~��[N�Tiү�߅�H�&;p�v��9�>Q� 5Eq������"P�Bq2�l���7{���c��={6��(zw(s,,�Q҂�N�s�������1%,ۿDh�޻g�Qt���Ō ��"��^<��}/+�����0�:���iQz	T��#Zϐ���c(��Hюqt��I�w�qFu�͘
�.�T�Կ����D������ƧQ��ѣ�� ��Q��g��/
6Г�����ww�����%���|�XL�X�摑,s��B(-˺u�ړX���3t.:�H��"��cQ���� ����'7������s	~�J,Y0�y��b[A���!����.��TR�Y�X)	&�`�"^Ҵ%�`��c�gL|޸��X��X��1��-�L���S����7���MOMѡ�K�24�����ex߅g��w���sI#$�����!��-�ڟ��kn�-*J狷��_��U�@�s
��)t�(�'q��kN�����/o������˻Q���?8�O_�\�M/mD�>�c_����v����5���}�p�7�Chǲ��y���+��4���H�K��
Y���/�63-�����_����� m~�����޻�����DfO	ڞ�Z�������c/��l��n����>x1N8�Pd�j*=���v�W߅׆���rH�
b�����a��*H���g(�R3dv�{�iq� ��3���Es���?n�3�.�:�Ht�"�d=��(~}��رu޵�p|��31@�eW�����:��ޏo{H���^��U�LXF���u�xh&����[�-��+�<�fS��-�ҹ�\&��R�-��;�jvP)Ϡ�n"'mb'����?!*�W陭�����m;��D3��}E,\2'�=l8�֮ |~O�i>��\��ϙ�<;����ޘ���(��Ή�U�3�v��lQ���l�&�鸪�;�������"�bP��<
���V��.���IC5�-}���T^?�\G��1�(W��D��n��<,1�Ѣ��ؕTbdX#@������K�~�N~��\�B��9!�9�S��u&\���yIڽp~�UJ
�%L.+�HQ�4���^r��<iB��tK��2W�D��@�Fk����1�`���Ϟ;ǡ N m��g[��i��r��iK�7��K��󦞀���&ց���34��1����+}3�\�ݻl��͠��	N��K����HZ-yj��MU�F�f�Y��Ѵ����+X�0l�Y���z�	]5��i���`�P%�G̜fu�4��y	��K7��G%%�)�~/�Sa�PݺK�lvV+�5����p�����'���%���fe��}*���N�}t�z�Y<��VLTHd�"�ΣP�SUyK��(
�vWI���H遪5����baR�mD0ȾV��*���h*��<Z'���R�n)-]o�pO�^��/ϼ�}{��Ab�9�ܫ� �S�>�0Z����;׻�mT�-��Ɏ�����7}�9>�~��Wh�cn+�Gu�hW��h)��RL�+�9P����m���})+A��5F�x��`O��gZ-�w��	���m ��`���?� �}�Z�;�`��7��b6���(�9�54��K;v�����ӛ_�ER}�KJ����L蘎��kiD�K��/L��A:�{���A�t�"�@`ib�V�	�5QV�?�p1F����B��H��D��K*�$v�2OO6N�F��\y�L���H�w�۰8�����me�h�^�~
}���S��f-g�@�i ��wvx:�i#W��Zz��L Zb�5���N}X)RY��)H�p�"�)G�(~�%��甽���h��b2�R�3�L�:5)���^* 1PT�#�af�������L<�y}E���Qc��Z����vS*�$�O�NԔ�A:�%��&�*�W��YRyuƔ9��#6>|F��u�3����R*�����`����֭czﳻ��+oĶݓ�4:�nﵑ���ulԧ��B�h�K��W;<2'ƺ�Km��j�����~ &Rr���,?8A�#�D �^,�5D�G��D'��N���vS�Z��)Ě8t�>\~�x�0��aa@hSH߯XOpn-&ޛ7��&����hvsh��r�JNW�x��o�B1�=�c�^�5{H&���WF�W�Ͻ�Se�������H�3�;�Gh��;��;�S] kZ�7߹��Њ�A'�E�0�$����ҙ$pG��A���Vݲ|B���k��4��a�0��|�O�{g�����{��ʜ���׎~]W��1|�_~�ݻF��w�a�����.Ú�K�3�
��s���m���������&�U`*A�:<rւ`a<T���jb����G"q
��_��X:�s�n>��|�K_G���'��S��|��)<��sسk�q .ڰ.Ɇ�{&��K��[�َo���t�Ѝ�`��f�b�{Sg�Lō�B�w\-���;�r�*]��w�W�"+�"p$J=_�bA�)��:�F�Z�2͘y^�H�*8����/W\�S�e�ɗF���^�m��#S���)�@:���#��g��N?��r�Q�6`��|?��:�vz.건P>H�WPhjo|�L.��)�ؤ��-^�X>'��<�Gz����L�cJ�#����dƔ���J��@k�h��)\�H���4`J�L�C�`�
k�e�(��W�u!���U��k_0gb*����E7������P8��UP���c�4�M#�Ni�3�
J��%?���j;�������d"B�fm;u锶Ik��eS�j+U#�y��.�SѸgeD�s����AU��ʨ�\�'2��j���Ȁ��:�KY�`���Tz�J�RTЄH�v�K�#�Kվ�{�2����TP�������i�M�cJ���(nA?��$��q�"!^�zI['M���~H��(Kr`��fJG�q���Kbvd^ρ����`��,�ӻQ�k�@H��w�0�}3�6�mUk� �c����uk��8�Φ����?�w�ԷF�;�݈��$6mۋZ;�^"�x:'��� �|�u4=�퓢H�P�t����
��@���ZXjv�m$ǌ�oX��tVFAo'���i"���^��w5�X)A�A����0�
������h�3��!�P0o�vP�2�ɀ�a��S����,� ��{aH��(�������k�P>�QK#�5�螒��Nݵ8���J��;ɺx*x��g�$�H�E��۾n���j3� ��ᘣV�3O�)������Pk^�`Gp��$�[�/�����xb�+�;�@'هF���	eLHNŸȮ���댓�~1���,{1���黾����g�x�}�s�� �i����D�jo'�TZ�[	�,�E#�ϒ�(7����b�&�h)*�\��s{ΓN�"�L���3"��\
�8���U�u�!2�o{%<ẳ�qu    IDAT�5�n��D#�c�y�`k���~6�9�x�}jA�FAn'�ڈp�ԟ{��̙�����"�	�3/��J�J�1�t19<����瘯�
H���N�)b��;�.�}�E.�|L�1mL���&�4�߇DI�)i���>�$��=��mB��F[��?�g`J��L]j�T�כ]\��0;��
L���A�M�),�V��.�{ݡ�v�������߃���fl�3�F/-?��@B�'����ڢ01�&��aiҥ��4 )X���]�+�&'+K
տ��.oԚ@y�����Uc�6+���	���+��.gf�D�<�%�q|�c��s޾F|��EE�����ؖ�F��koy���P�:�!�m����r��V�*��6���)���W���}ҁ"0ݼm�������;�5��C2������5�h5&�j�����_��$��^{����ނfl�X�b?���1	wI��a�4��Y+C�#��
����֫Sh�!��W��\|�*�<zQ����m-��
��W]{+�����Ƿ��ylX��we~���p�Û�F�� �)H�A(jb�Ff@B�G���1Q'YI�jRL��`L�*���p�;��z.�4d�:���{_�֕ҡ$�u��;mL���n�ȃ���x�=�B��ё�M;{���6m��IS�5�y����������Ӑ%��dcۼ#����T�����L �At��s��FQ�z�
��i�TC�5�_�}�Oć�9/�'^������՝�H������ߏc�>G� �:��0�&'�|nz�14*38댷���++~�=�'�m��w<�j|>Z�<�������H`"�7�l�::��Դ�d�%.]�^��X�P���]ƽ�3*.;V�
ZӨN��I3P�@��G7����V~��.�Z�=�R��cJ;���'R�9��ah�sK���!�<3Ö*�y�ԝ�*�:K�D'<�9(�t�(��g�6��RqVF�Z�Je��C�j\�^8�p����!8e�OA)��JQ"��4u6��T.R���'�i0�Ѕ�����g@Y��ͯ���vG挂��uI�U���7-�hE�E%�B�_��y\��J��0D踶|vl���<
���)��{­N��������4���p�����ܓџO������COo�d-�XzZ���ՒG>��	��x�3B�v��*5�g�AR �Y.�.�%���d�����S�(&V!�R�Y��,�ل�S,�Q?���h��i���r.���p��sE��I����(�u�����ԁ�;���qյw��L7QD2ׇL��L�t�tZ:����.g��KG�h�A�� ����))�ٌ�������Oj�n�b��#�W��҅t�j�:�Aޥ+��w�R)�e�;4����)�(��F�3@�,o�3�
��;�o�E/�UݓRz��)��;{v}٧Ӄ(�<�56�(�#���=��5����<?	 �WWl/�~�+�j3�g�E�G�ZH�v�O�.f�f��z�A�1�L����w�u���j�<�ܿ��}�aEEǘ��+������=�`���/i���|��,��=���-�ޕx�G�6`d|���<(�5�EL�O@ʴ�W_� ���s�kf�;�fj��{��I�)��9�V�:P$��Kfe�� U����?�g�}�\\�ߣ��{w��>�Z���vV��л��a��bio�Ⱦ/����Xw����%���b�,��Q/˩��i!	��̱}މ%�r>�b��*��Ǥ�/���t<���65��,.���/���*.�u�.�Y�N�tʨ�]��N�E��T�T_	I��R�gB��cn�[uџϢ����>U�ϟ�e�.��N��\�fL���=IPW��g�W�)\��v�������ù'����������gv៯�����N�jw�hw�9�".�a
e:�-ɍTt��!��Dɖii������-���h�r�uX];t���A&�"�2��c��F�"�2�g�ji������!#�Q}(�N�e�M�Q�5�7�X�a�F;��J�wN��?)ղlab��T��$�a�*/�F�"^���^�ɖ����2��6jd�����=��u/ʭ���]� ���FC{�@��W|�Oq��ʅOPt��/�
vLs�8�J2�(�"&�6���TcR����yDi,�/�E���VF��h���g,���8��hN�W���&�Ͽ݀_�q�>~٥���׉E�r�͢��?��.<��Z�A$3�����|�����������N�P�������N���;�h|��caI�*-�o�~=���_ �#S��EQ��Qo���Y���}�p�ʄ �
g�c�$��j�5���o
�u�JR�P�ۯ6C*������~��c���N�&d�*MOJ	��_� �3�:���̘\�z5��6�h7;h�Y���q��$�9x.~��S�����}�
����-?����#ÒKP,&13�NZ�+���3O?��n���:��ذ�$\~�{�_�+)0Az������x��t�8�$1�Cg�"ѣGW7 ��1�it��}���M����J\���ްq�Y ��i���gʲ�ż�\$�
�U+$	��+ŏL{�T*"~�zCL�`�Z��|�����^��`�IRZit~'���s��|j�T��P(G�uw����K�N ΂D�(���^�N�{����ϗ���-�`��h�A`����G_�f�x��5I��ܭL�rM���=!�:HhC� ���Ld0�as�Kb�ɋw�X2k��Ph����u��!ڭ	�
M�I0m)]S����s��??��|js�q|�����v��*��������h�����Ӌ#͎| ���ڳ3N��F���ݙw�dM!8RW��By�6!�:+�@���!�����=N�����N�ic�do��P`c
����&6�m-.8g=V��y�x���E;)���������_=�ۈWw�Ҋ#��C:���\^��q
�Q)@,�7�~B:h6���zr�)��
 �x�,`��K跣�(�o��ߞI04� Z�uf�a�G������l6��
�6�T\P�	���!w��X�L��Y,	KZ�>J��?�]XU�V�}�JC�y�����0�]k�Ne�˃� ؤQܨ��vxn7$��ے$�#/��i�LOIA�'8kanG�N;'w�.��^�3�/t��#��%�����^��0m��D=�f<�X:���ɬ�#D��	He�T
���9Պ�S����һ�^X��'@�5t���	�}7w@k��$�T���[�H�)uM��eis$��i�Hh)���42^�L��:q
;)cFf���(!��j�ǩ��&��hE��;�����>��#���n�ί��^��,ϊ� f��Z�����Y52�d������ލ� 9���B�&}��nK�\|Ɣ�P|L)�I�̝�DJ�$�3i�k݁�0�H�%C���6D[���\���t>h����Tǧ�Q׍Ǒ�����|�Y�[��.��Y��v�����j�U9�\�Y���`-x	�WسI+ �OI*/-c��,"��.�tQ��/~�<�}�6������'�75�1������������~�\ɗWdL�nm��[�Ψp����#��<�6�-3 F-� xK:�Z���OpS�A���Hu�(w2�c�P��A��e�^C�j��	\|�q��?9��i��Ö�q��
7o�t�-�k��L�Jh�Ҩ����jcx��f'�L�O:���_�Cu52�Θ���!��Ͼ��]e����ݓ��W�'_�D���˗c�;���u'ct���o��6?���̇��g���B����m��o\�fb.��2ْ��rF10дu�J�$ef�����b|���V)�^C�=��|�Cx�9�:0?%iYo�5�|����9��{�5���ކ���Z�9r5>t��0�_i^n$��Pn�n�/�ۈ�7���2��j�.[&�s�������4�4�tMc���!�_��yL{��b���]���W�ŊHf���Qcw_TJ�8e�A��G>����CFq~0s������<���O��{6b��B:_J�����y̮���,xB��]�Ek1�pGPJ�.���@B�~���'�f���e�LϠ\�Iu�獀C�:5t��8�~�����LeKr84��M����>�uo[���/�}��V����s�xm�.���x湍hT�x�����3�!�2j��?2���W�e�u���Ԃ3EU��K*-����	ԦfdR�_�iF��?�+��U�kON��E�wl
�Z]b �i|��T?�h��EL�:�V|��4F'd�T�����I�UgM�P�\�7HB��%v.��(�#[��	��5�~m�j��S�ϴ3�ϖ.��:�X�\4�I3�v��(J�,j�HǪ����b�E�'U�ul���p�Tb��H��z��,�e��}�:�R�������PK%;J�r^K�#v-�eJ�:��IK��&ɴyd���&�O<y�DF��VΥ�t55�Q7ҭ�0ؐ�m
�0?�+>�!���rc����[*�ꖇ��潨�dԾ�~�&����Z��f�M鞊���T�\mg�R����;`�+$��� _�(�:z��X������]/"[���v~�R�m�׬�S�B�5�Es�8����'㰕�(2ސ�O��
�� �e`��I<�؋��'�s��Z;$K"����M���E���T>�-���x��첃/_� F��A ^���]`��̖��;��ܡ&~���Gi��n�]�F�g5ٵ؃x/���uf�rq��Z
���ޙ�������e����<��{	|w# �_ԁ��S�(E�+�+U��֞�Q+�E�;�N���hh�}�u���Y�4�U)����R�%e�������9�8kV���	�R��o� ��9��6��oUq�Oᑧ��=�h��h�2h����5' Լ�ۦ�vc���(�Fz�^`:�Ju��[�L��lB<^D����Zg3�K�﯀f-{�*��I|�����fK�Q�0�e�8�p�;Oӌ��I��؋oa�Ic:&jl�Ȟh<H\�e1�k�����Wh�w��=�h��?��Q������ZX@���rPXϱ8iQT�Ƃ.��Q+*�N>���ސ�(�}Wa��σ��)3�E�E�ꖊ�&�n�c*�"�d��PL%�c�lcrH;�\Ov73}Hҁ��e;����q)S�1�t0=2����Z�G���K���[ň2RDdV��Ҿ\VTy���Ɋ@S��R	�� Î��HÄͥ`l��/�-a��c�hNbI��/}�=��!�O��c�)u?��+��-�b�d�̀��b#[HL�U^�]�`Qs�I0�����A��,�sA��H9SE>{���Π
���qI��b����>�YT��s�(#h�9�K�s
>v�:��)0�����/�����?�ͯ��I���![ ��* ��C���G�"=)��j�Y�|}��+:�yi"�]A����/_�I���3S�J���x
��q?F�j8���pںc1wa�'�_u#vn߂���pĊ~9Ȥ�<��^|�Wc�Уwd*/�	V`x�}F��v?4V1�j��2�nL��։)�Q�E�=��������#&��lzW]+�"��}���Us��x��kp������!.�*�*L%A�>dV8�rx�M�����ߒ�<79�H�p_��vl�*�]&�d:O��(T�.AE��`ʎ�.gL���a��7~�z;%jƙ|Z���	y�l1N=�p�z�AX�l.���*��|Ry���xu��o]��_�D���X��S� wY�f����'��p�QiD	� )�M#E��dRh��	c��M��0�33�V�h��9Рإ�(k��i��������/�<:�X��.��L�Zs���3�Xx(��ر��X��}i4:�+o���g�C_!�S�[����9|?�~�˗q��a��C'M�͔d��fKY3e`" ����>]����C�R��%S�Q��IѢD�����E��I��
L��ȧ�cJ��N���SyY�P�!_�W��>:.4oI&�J�v0�3���"Ve�A|K������E
��^��,-�?U���Y�WlaXȡ�}J�H�蒪f>�
^4i�Y�iV�niv�yv��Yo�Li�e�k��b��Ku��vVC�������E��:iQ��W�eߚg��g�>S�	�Ϙ{��H����ˤa�D��9\�@B���doa�J�[ޙ$��� M	��E0m�kL`������q� -��k�.�_|��u����_�t�l�輼o�����̍�w�v����:»����kx	����G��7��5Ѯ �ꜩgUg%�ZZVȭ��	L��g�� �1%~�G�g�v,�^V,��=�j�Qq�nO�($Si /�Z�s�������M[wc�ʙ�lБa����h:pdG�2"�ƛ�����Gp��5�A �[�k$����������p]���M{Q)J �^'�:V���$��?��?-@p�bcx��tV�əM�7��]���"3�Jr�m}�m�B�_O���vrAB�Rj/4h��3�ӽj3���0�K,���h� F	��q|�J��q����$5��UG�6��bkV��O9��[��K�ȧUiWWT�A� :������g���G7b��!�W�6�9�<�قX�Œ�Ԯ��W�~)(D �>>]����C\���S�9�GN�f�&���{��3"0�h\}o�'v`*�X��&��T��M��=(��Xw�A��ߍ#�#m3�ަ�O�~'^�xe�:/	���0W����S/<x1�?���Pl��Vİ/ ���}?�ߛ�;����@�S�����}!��� ��כ8������X�
���=��z����f[��)�Y����KQK}��8�
�K�Y$-L0U]���/Ȍi�T^������tQH�)]f�86UF��?���}0=2�,?��E���|�z�{Gј�JJ��r�4� Y�1�gm�V&t-uH��c�⸀�v����`J��u�ل�n{o�ch���"�d�R�L&�@�GYx&�	3�f��s5j�B��B�`0�dA�ö�+���$Q�F5y��D �Q�dQL��;HL�c�I��f?�էޏU����8������kp����d�&����YĒ����Җa.���y�b�ըt2-���#"�cC����WƅV�Z�龭.ʵ&:�8��4(�ų�c���~��q0�>t?����������-w>�^b�ɒ\Ĭ,��䳋*V��۠�N*�@zI��Ԯ�ժ�L� �+���>�v�w��}�z����@<�#[�?���jiYn����8d�
�8m�H>�g�<��Y�^�ꦧp�/��(�ꘘC�:����B)�͘DZ�3�F���U�T�zu4+Cx�ۏ�?r�%l��O�8����_at������?
�-��t;�؃M[^î]����hn�u޹�T�>p��y�������/|u�9"�AO[�TJ�(��[���[�{�"��i1��f�ͦ���N�I�"+�>���b��g�I�m�(Rr��&������1���?_�q�,){^�`�E1��	0�`��!,_�}����hr֌3Ze���yo_������>4�)$I��.)�B�Up/�ttM>wz���_��|M�!SO��V�%���}����Z�g��7�#�j�2M��Rշ�.���P�r1;�<;j[\�F��n��?��3:���IiEAW�*�rQ����������M�A?�Lvh}*
y�y!$�ce�Ί��Zk�K|��Y�Ƅ���GOۆt��Z㊶n#�v(���jv�\y�7� Z���;�ڡqJ����C�Ω<��M�T6��8Ieq����_��p���þ7>��m��c�ʷ�����iso�?�M�Y�KuՂ��S��+��r�I������]�������]mF%d��d��D|���)xR�����.ډV�,��ĥ��'�Dڅ�� ~�N���g��JRk�m3�,N,a���ք�Ž��2�`*ϓ�*�{    IDATG�-�fdd&ўƁ��O��|���՘S�B0�.�y+�x��b3�F&���߉�q�߲㕘̑Q�)P�4�d6��fL���R�-�� {юSH��dtnRC�NnkE>V4�u[�ݹ��{��;�bh0��w��x��T�b��,�A��X��8f ��c�E�a ��(�ɐ5��+^���R��1�9�������������|�MYv|d���o[�*;���p��r�X���*ˠ�<�L��q΀��e2X�z9�y�8~�AX2')R5^�R����w+4V$�~n~���xy�읨#Y�/~�d�v�T	vK�|�X�z���zr&Yx-���X�ϒz�`�l,��=��ʹ�Xt�.���=�x�:
�43���3M�ƝN�%���Yn�טF�9�����/yY�����לS� �+C�7~t{~'z�~ētV��uʸSW
��|(M�`K0!0c����d��uM�����y�N��j_�� ��W�&[���1���*諈��ِ>�*�Vx��?dW��p�ђ�Eq��vL%ס~�) K���i_:�t[gD)�=@�a�TD�/�v��T��\�&fWH&0���.��jST�[J��Q/�*o�]&��"���r��R��Cs�&8�q7O�L
]�Q�z;Z(q�Y��Ryɪ�>Aj��@�3�E����qƱ+�g�#vL)�s��q�ݏag%�F�{-��U��qH��%3�0��"D�<��/����3�G�$��J���
��R,�Q_K�@i��D߁L`Kc�<��3��ܞ��b����xφ�1�S�{���`�W���]�RZ�D��ȱ*Uʃ�����xc��=V�,�pʁ��Z%\x�	G���c��m�B�"���R*vl���xuw��x���
���7�M5|ퟮŮ�6�� 2@Ϳ���c T5G�@����9��&tA�[:,"�sl�F�:�d������_�Rsql}}����s�����y�
����p������8��UX��$�0X�UX�����#�շ<���ގ&r�řlh�T���[l�r�=�2�9�Ap��f}�� _���a�¤ #~�j��׏chd'�r2V��� |���	��܌�=�,f&�e&eN!�?��|�߃����)TWݶ����h��dR9
$%ys; ��l��D�ɏ^^�F�	JS��s��ҽ��@�+�jU*nR��� =S���ʞ�_�m�֐O�qᆵ������H�I�R�����M���+;p��S�rq^������#�Q��&�7'�_=���������з-��a�Co,��\ 0G�\�ϙ�1�d�ˢ!v1.p��cǔA��P�2�㤚Ӫ�'����	1�&�WEy�Z1j��~���1����$ՃX�i�M���m$���A��f��D�.@Y�U3�ƨ �%�" a�{�r�1�e�R�]>��A�1
m��Z�St㼰(\��e��.��z̥`g� z��ɡ$�F�b!B;z�{W@b�	���;P솹Կu,I	&#F���	�y��/jɖ�)���Lй���ɲV��ʛ�\�R޴��P�,1⠁ܮ	�H�cgT:�2&�E�QA�S�`����$\v񱠶��NK'.��M&Ăj�n�'7=�_޿Qf�, �Ϋ��PR]U�~�����d`J���٨���"�"ui��w�v�$,�O{��q��l8$ka��.Yq+ |B�	Ҏ$q�}͙a��[8���x�����5�`>�>S�0/g���5��z�3��(�ß��wb��C��t]�
�2�l.�� ",��xF�0����'����gEMq����ۆ��HA�^4F(���޽5��-�X~�ig	Zs+ �>�������{�4 4���1�>�W+�*��jк�#�� ��%2�3�F�As L�tM"1R����w�\��*��h��=`�8P�LaMi��i��]�J�.G����j��~�!�q��������Z�
eT���r�O������;ă�lD��y�$s�Nd 2�b���;���*q|ƨ�zV�Z�����&������r3�І�wu%5�+e6�OV�V�P]WJ�Ҽۭ���sm��>3=�T��R��w���x=Y�FN�a�߶���Q�'��[-|��w�闆���&R�I�{E�=�q�\���̬�e�]E���=K�(^pQ2W:Q�� ��A��7�d��[cC�(�l���2�³�k�5���=�rV��eςtV�qH��i�|L�ܐ�M��R�.&��f�TD6���@ b��7 ��1�LrYĚuT&&И��VoJ�U��}�dXv�`����:"~ԟ�ɸ�tLgjrPh��S�tI�vU^_++V��2�����IB`ڕ\$�k ٞ��B���ǭ|�ܐ��W��������/����F�$��x�� :K�j/�RaSɆV⼫�m�
ۻV���1��px_7�S�t3�Q����Y����z��3���UvM�H���.���}�Z,����Z�Ҫ��L� 
�wC� ���o¯�	�VqSH�����fie���Wf�ʈu'1���w��(����X� ��B���:�\1�$>�iv���;��
��&��������nB7�'F�|���a~v�����:���S�ZH_�ں�2��B���N>�0���]xy��$22��h�&�b
��
�tZX�t!X��[Zml��ɦTwx��M�.ㅭo���B�u=�z���*�.�R���АZ�S'Q�:��g�ܷ(�i&�ݞ[K��b/%RRI���?\�G�~	�Z�T��28�؃����߯ kC����-~q��ht�%Hf�H�2�<[o�,	bN�u*�%ќO���R�,����v�#�/�jE���Q�Q�/�|h��w�mKN%=v��#XP.:�T�����iJ:NS��#E���-<�����_�3։��94"9?���U�G7=��ވ���("�+!���'4�KW�;�n#��HǴ]ֹ�L���%�dƔ��B]:tZɔBA(���jǔ�>���A�I��j�Ne景Rm�S���[�H'�ڡN����TF�[��1P����k록oM���2k�?���Y�v��i�����W���=��Y隒�(���"򵢲K1:�s�I��ˀ�V�fKD8c��q�kUY;o�;�a�X#F�1����:8�E��%��Ջ͙�ϐ>��o0�������j0��JY2Kd}K��H z.(�N,�کR �ɱ�K�3�g'�[A�T�m~V;�:���)��:i��$Y1'�O^r6�8~%�L~M�Á�tN�~�����p�=ϡP�TN�)@ŇXi��H�R�r��G����O��麩=�%���:���>{]�pDBi��ZR��ڵ���J�U�ឧ��l����06��tj��7��|~�8u.<g=Z1(
�,
�0���OÙ)�������R|~r3�~qv���c��*Y$�B,-��ʼ�\(?A� ?�w����\���*������K�	�w����l{9�k��:c&�]�9����Q������P�LJ�N+�F�V԰ן������i�|=!�1Єs�+��~�"�[��{82��aK�\��6:�3�W����GVd\�ñ,mk�I����3X:?���w�u*�:l%��O �څ<�ݾ�M|Z
]Zx�{~���y<��F��{�V�L	�lI�b)�i��� �-1qJ��l>Y>�%.6�.�f�fP���h�W��l��Gؼ��w���X`�5j�K.{D��ļY�����"�	9�!ֆ�1�����p|�����e	�g� Z�>��^|�'wa�X�v�lAĢt�XG��l�@�d�\�	�.�M���Ht���ұ
t�J��vƥJp�md�)��,�1��=���f�ܭO�����V�Rb�S�5p�3 Օů����hN�E혒�!����:.$b($(~�ER:�èNNJ��ti
'�Jy(0U��>����c��ч�&��ZS���IM��.�"���ю'�t�E����B%�JU;�3�W�H���*p.#3�m�;u�V�ҙ}��إ�uQ`JJe�[��?~!N?vy���,�{����j��'w>�k�~C�tL)��J���(]�&����+V﵋jۅ�e�1�%QQ栚ii��9zi�}��M�,C��\S�6�F�D���l�^hב�U0�i��N�{�?K(8e�����#�7vE������[�����K�����P3Y���j��d��~��Zy7J��Xw�w�98��w��E��Y����������gb�҂�H�̜o�jh�w?��><��k�&K�g�Tg1�ζ���Th���s�Z���趐I�Q��0U���M̊`<�FK�;ͺP�Ę�G.��6⽖̴�O�Ǔ��YB�����!�) A�*�K�E���jh�+\����4�-��k��G�zE߾�ϰ�Ī�Q��rЮ1�w�C#<������k��F�)	+��!�������뗋l�|쯮���g����IJ�~�,	�g�.��H��8���i�BY
{�q5-_�5^-���UG��F#��J��j��/0ծŠ����T'��7p�Q+q�9�qܚe�+�gJ��m����;��O����i��]0X��o?�OZ�e��@|ķSoc�-���p�]�b��C7;�T�<�29$�9��:�U��J��Q��B}lB��m:_@���|QݒHM$�$�6���i�T��]kȖHH�@��$�Z诞tJw�j�Z�i����H)&0U^έy�٭����,+�Hbޓs�`G�݁�e�Δ�W���:��1���s����X/���R~�+�27�IQ ~�� ��H��b'�h3�FC)�M�b��4�lGi��6[|uJ�^�~ٛ�b��j�5��F]�����'�A��(����W�_M��������qS_��C�O�@M���U��kW�%���@��0��ͤRB�oq��]E�5�U�O_��XO:�)��Q����������{�Ƕa��C�8�g�RH�Whْ7�@�I��& �LT�h)kg���u��$����M�
�bA$׳�T�ٝ"�̪�R�� �d���,�]�^�4V� 睵�>s���{�/�׎ε:X��P=��N[^��o}?��'Z�u��%sBq�ˋg�wr"��X���w��9�U^Ψ��νЩE=��wStG:}ovƤř��i�f�/l+�ȼ�t<��$���L}?p��h�MsK�f�|F�!�T|K�3o�:
b��Z��`��EjXpR�j-���΢�O$�����:�B߷�e�@k��@��z]��X�i�SZ�x�sj�V.Ć��S�?����ǑSgM���zW^v*�O�ב6���p���bӶ=��H��!��eQ"��]�]�4q���~	��>�+�K������X����8� T��u;��c�����^*=>��� �B؆f�;PF�\�~�Uԫ�hUƑ�Uqґ+��.�)k�`P*���<�=`������ݏlC#֏f��N]	=;�b��		��`w��a�X�4
�]��=�������'HqN�V�&����@`�9z�<��/"�Ж����%e���gX�������f�EÅ9��q�y��a�^�"��"��]��I�П�!��`r�^��RC"�D�T�9�d�1�	�R�#����l�z�)�JMQ�`Z"���,��j��f���:�P@�\��Ш��
�7��#S�(rű"f'����2�8��c�d��G�:�I,.4��O\�ӏYtL�[`Z�u{��۞���<�=�,ɢ(yj�X���_� `]S�{�K�T{3�v��>=��6�ST��:�KӒE�M��ݥ� Z��yS�Q��錌�û���&ڵq�m,YP��kVc��a��1�'b����8fjml�1�g_|�>��҅i	�mtѾ���x�v;4�S��G��T�K��l�|�b)�,Z(Ԑ��1��Mbhl;���P,b�~��r�;ЏR�$^�3�F&[xc�8*��9v�5��9R?x|��߭% A�YI��#ɘTՖ��B~��,��J� ��{ŝɻ��-�R�K(3�Be��zRԍ����6���G�J�Zݗ�n��B��̼�=5�e:��`24��]���0�ƓTrh_�B%"��^�����_@����"�N`�¹Ƞ���{�u����Ol��?]uv�e垳�ِ[/�\|��� g�CQPS�R
U��TT�ia��jx�:��|�hho4,�����L��[��b� ����(ڍ1l�/e�`����1�T[`9�49�^$ͩ�@�UA&�C!G�ԾnuZ� �F�@���\��9���	�� ZlX��畑�^���ǛMT���6`���ѿx���1������_}�]��JMT}[?�|L�$�T:�q
��ޞy5��cJa�n����$�LjM`j���K��(���vDI�b��BH�-}�@/$ݧR��\��Q"*������N�CS�H����Ȃ��G#��1�L�I��]��u�%ڜ��Nq�:�V�%)p�x�Z��Y/R�������0X��wL|n��>U�O�s.~��d�߻6��EtzjJ��3X �;/P�<�I�{b�ʬ������H~�?�(}޴�"!�H}"e�6�^y7����'?t�^w������+�#8}m��Ϳí�<�r��xII	L���@I��`Y ���!�~�4z�8DV��\��,��C��<�+�	�
:iȤD�b�l_Kbh�;��^��V��wq��$Z�1${�d ���3q��c�xnF�	����p�+dIb܃1�z�%�������0&+�� ��0aN@?���,���Ȼ="6��	wM�P�����H��ɮ�=���2c�g�a�.tt��<�[���;�Rd�N�%ݚCX�d1�z�����(F����ޜ�Y��J�a��
�� ��T ��Ě͢��M@R����cT�^�5��~BTI�d��s�L�x�zjvE�B��Rf�re�6-3����X}�R�8�pЊJ9�_6&w��
4O���:,�����G���=��2h�����bHm��Ui7��E,�;�2�0���S�>_�Խ�tj�9���Tc���=i�Z!��T^�i���EOߵ����h���I����c�V]�(��{�OTqֺ���?:GЇB��o$O�`������q��[1VMQ��XF�Bm�¢�Q}[���y���P/tw̾� �k�KG34&+a�r.g.I�⑟#[����ʎ1��zA��G.�c�;ׄ&	v��F�R�1�ٱ0�kuT�3E��bX����u�����P̤0��V��Jד�T�q���b�tq����� ��S�����>���Dx` �TJ�8|��Y���y����<�A�LSN陋/dT�S�~Oj<�=�����h�T��W��K}�q�2�˙�w��.�T�+�n��i�nfPKrƔM��
�f�=�	F���H^�9�h`�c>GK��*�'��Z��9��<�[���ͅ�O�BL��d�T�G�T&�k�!Acf��J$d�9$3Y:`�R�c��C,YD<UD*��PH�ڃ�#�66�;Bujw8\^G�d^Ԥ�t[r����9�O�k��҅�=GyfJ�+��h3sO�+�P@�M�<���!�J�~x� ��Y&}[hUM+�6�i^W�?�j��M,����Px�=�V��}IҐ#�p��g���k)y�s�
K
�y�a`��Fc����,��C�{'N?e-��RPL����w/���=�[^E���D��$��\�n�������l!�����&Ff8��E&[|z	�d]�d�}�.���ɧ�gJ���$N��'M���������]p�iX�P�+&������%���u��n4j���&�Ո�����������LF�;+ԭ�E��%괚�e�?[��yȖ�Kf�e���Z��$�փ.��4���(��e	�옒��I�2Q`'�}v~F[z�R��2<�.׊T྾�c��k�F��"��N
�)�t��&�iSUť�g�4�    IDAT/v� ��v������ׇ�)���s
�FK=\����l�"jI��N&f�$R��;�3//�������ha���_�b�	�6(�K��MTī�A�Z��q��GE}0]���  ���w�<�(8��fx����[t�O��	�ȩ��%�4���+�z��v	��Tۅ:���SE6�*�#^�����`{^V$��#�ĚS@e+�%�?q)�~�J���3�~Zvh���L���?�����TY�xS(�
o��.���ܕNI����9d����	�H�,R��0�j��y��X�ɶ�Iy���
�ݖ'L
#�uS��l.绩ދ.G�Ѯ�#ў��W��3N�	G������u
��:�m��D���n�:x�q<��lپ;v��t�-�e�gEԃ��L�X|bl���2��g)1G-Ǣw���e-q�����^x��ߠ~�$�\Dp�ї��a+E�z~tk���������I�.�����|k��bK�[iBߥ��X���k�AT�%��i�Ħ�X�� ��v�-ԝ���>�/���n3cg��K��j k�THa��8`�b�\� 'w���|*�L��o�H*@��l�R4��[����3[0^�KɌ:0HQ6�)���"�� ; �"V�>3��a`1�#>�+�{d��Ne���<�?�i��6����h9;p�G��+�Yj'&���4I�2��8����ǿ&V.�K����V�?��;v���������A�2��g�ă^rC�6?m��Z4	=*�;�G��h��"��E¨����`tf%����d<�Fo<'���FZ�Ʊ3&�̺ϓ,zUT�_�L�`����k�qʲ ?��GI'TG\LYpN��J2 �J��K3��|:��|�F㻇И��K���~�̗j��6W���XK`J�X���Ĥ��5�rO�rH(��9�|]�&^1�E_.�v����hV�rg�YW짢0=�Ct���j��Ɣ�m�'vzp�6�.&�P�����E8�eҙ�ΘVz�^1��WO��{���N�x> ��u$�Y�JI���X����������9�����J=�A��:M���Y���a�kN���\!�)�
.k�8���F�B腤74�z
�5���*��~L�6�E/F�*RX�����q�'���s
��3��vz-�;MI���::��4A�L�`� ��
���=MMN�IsI�r%�0�ΣP�@�{#���g�n�T�D`� I��A��J.��Z�o$��j�]�6X��eHm
�l��S��j��.���>���]ڰ����^�:嗭'���f���eN<���)t[�(ezX2��#��� �U�ؽw���cSM�P@�0-����0��w�+����t��r�ꛤBP	9-s�ywZ��5`�C̞ؒP���T�`���A��@�^1 O��oL�m-T$�(R�`Ze҃xP��DE/1�xw;N9�*��t��R��w")���:萀�[��^�!gF����XD�0XR�k{���CvlmxU(S��KEp�����;��q�����Օ���{����9���Y�$ �F��vၲ�\v�Q�TttWT��������.�-��6`ƶ@fFB�Y)4���;�k�s^�n*Z��|����=������k������N SVL�P�`�G�_��8S��Ǌ�u�?��b��b��h�
����)�u�!�Z΃��[>.�.õ0wTO-�W=d����8;#���;*v�b����̻��i*u�[M�M%A�����yrxI�L`��ꊹ\?��,&�	��$�$W����RK%;~0�LT3����Lf�D9���IĠ+c<��ܡH�=.E�l�x�4-�.Έ`�I:�Q�U5��tz8���w�t"R��I�K��n��H�EO��4H�_6���l)�䨿@e>E��`>���x7_�o����u�:,pj��?����������W��-lM:h���ȯz�?e}���S�[���|$*�z�ѵa����w�=��v���1���h�'ɼ��O��.�h�� �K��]�|�	='��t��\gk���9�l�� ��^u�Q��-��[�p;.۟�5�0#.�������0�1I��)A�8{q��^:��=�>��o����?���N�vw�{�;R��-	C���;���Z���=*犅�f�y��t$!F�$�n�X�Ȟ��� R�4���Iy3\!<(a�e�D�ftfzˀ7���g6�� t�;�� ]ڬn����ʵ���a��Uݳ�P�3�g���l���f�.x�MF��vP�ΐ�&ؿ��[_u5���;qݕ��+���+m��b*If[�^�����$�Xab�tc�ڃO�_�y��ۜ`VmKU��%�%��t�.TO@m䕵�؛L&o�Xi�ݪ�qOC�f��b�l0����r�]���g��EE:� �t�ZsŅ���g݌'��9罏�h�� �����{�pl��.\��j�"(��3[���Ǘ|�Y��$;���\�{�c3R-�wC+]wTN�2F-o�:*HK�{$�ag��I�h��a�%i�V���(��宆+�/ҩ8]��BY������<�M# M1qɓ�c���U3�e�9��m6T5UŔ�'�)�"0mT�b:��������75�b*`Jh�{���R`,Mʛ��� 0���	�K��u:L�P�:�$�I�m��v+�á*������4��ǕE���S�gr�sȌ��j&�D���pp6�6�-iO��O�?��}��m�������I̻3�7909�r^����~1����R#�n���]!OT���.>�n_QU��¥4�)p���>ɥKX�J�C��OV�ރh����A�Q�9�M�&��X����iM�%m~?��\����,�<��l�ă?��t��w��ôp�[#��$s�$���c E �7��<,t�Pg71����*{�/>.&������O��.�R��`zS��`���L6����%8����x?@����@���:X];�?�E�( 4�3\�Sv:A�QC�YC�һ��+�[f�P�TUH�%���rc���%�$c<Q$)A6��2�pd��Kx1��ɋ���d�%0L��K�J)I�`�yPٻ;�h)�v9�O�,���ùџuR���R��u��)W7tq��LQXy�q����:��zF|��&�K9C���6_�b�UP�PT��3��d���Z5)�t�ޙ�b��]�1]6s̀�����ǔ�(��nlaF�3I�.]y�T��W5��*�.]ҡ"q[C`:!0Mt_	L)�M*�m-�>&�,��Eeܳ.�:i�n`t�Lџ���|�t2�U�����4�9ݩ#Q���R��<H.�g�{��E#����	�s��!�ū#|_d����VO�KI��-�/?���&��#�i�|�Ő���Iɩ��v>�Ȓ ��!���^]���'��k���'y�֧��{E=�Iɴ�8?��r�#����8�bޢɃ}\��KÙx1��ܬ�G�x��&n<��?����ͯ�m�S��P�f�zOo �}�a|�Ͽ��i[-�Z�n�F.�#,m���$�
��A0��י�g����H<'J�(H��d_������G��-|<��vo�!��x+�P�"���t:&q�Gu��x�4V�S�t�a��Mw��o�G55_9L�e^|%�Qw;��"�)p�<��3��/}���8{a[ uY�e�Wop���f�#�ɼI��I�,�t3��\��23�L�����}ׇ9������٪�6�>3U���1�������h��9o䟻_��*ͤ\�z���*�>�A@��. �KQ��10fy��~�8���9�wUw�����h&�|�	(�%�d�ƪ�.��FI�c4ks�x�q������{��-7Á�@�%��9I�G��T�:�q��h�5��� �����gNb��1ES8��{���t�%h=ٚV^�e9����*�n���~O��8`U�]$����Ş���ܤ�E+��~ dϩ,������Q�buzs�f�>����u\u��_�����|�m8�Ǧ?p}��H:q�0�"yr��?߇'_�Fo�@�J*)k+��К��~��R/Z3f�1(�^0�(�*冩������Ek���[���ϋ��+�v4�H=S'V��]��\E�4���X�n��G�����/T�t���*�V1%�X�l��Ns�R)��jݩ:�D��a��Du8���&�QE��ҡ�7ØK��+_���+Y]易	z��2Hd�i�.L�9����0m��Nۤ�́)]y;��	
�y�L1"@�x���]\�M�jJB�μ���P�p\���?y�����C\y]���o��[ŔR^��dj��U�J������]PE��%�O0cG�rKL@��[�!��oA��!��@�e&�w�5U�lUh�C�����L�cJ\&J����,��Uv��fS��fP��Q���3�ԨK
��B;��O���X6J��Q3�  t��0�dpd��$�M�`�d�!� ��Oߕ�������df.ot��(�}Ș����OI`%*��X�9�U9��p2>ܸ`�w�U���Ϊ�QO�9�._bŌr�۔[��<ǡ}{�yq�O����)�䍗̓@4���H�J�C�����dfU%���� s��#�Y�����*�q�7ԣ�H}��{���$����	��s	mB$�,��6�U[	\j5��Ij�u#�1�-i�D2 �֭;p{ŝ�i2���Q���JA*���&8�t��#�U|��G�RE���}�ϩ�例����3��67��W2?b��`�����t�0����bJ)� �K�7�H�Ã�ϟ�Fe2EC#V�G���m��Eu�%��H�+��Wwm?فjQ�*I�|r�d0LuT�M�$ �ڱ�D4@��G�1��FȜ�$����J�\NiɌ'�>n@k�4Z̩~���(��@�*�HR#)������>|��U�Sx�\|7��{d��$��+;��{��q�I[�@�}zb�����{�H�c�(�	�p����,����MTr��h�F�5�b�	�.�@k����{�q;:t�-�SU�(E��P����w>�7x�mT���6Z謬��6�^�q)�J:E�$�5b+�ݷB������ ���D ��O�ͥف�ml3��]�^�\�xc�X1/��L�z�B�`rm�/����B�S:��h��|���x�����7߉7��U�����p�n�@ 3�B[~1���n�&m�p.���������'ױ�5Ҏ�	d�7�Bc�uP��dbX7pJBRce 5"�� Om,��u�(�R�i78U$����⽐Y��'ܾ�-��%�	�ۤ8s��Y���+�𤕿�|(�W��QH�����?�cX"�R����F#���툉�x8�X`�$�w*�=�Q�>l5*8������m�\��^�J�|��8|��n�@�s�)&� �߃ּ��I��/������A|�k����vFT��A�ٖd�.��
�A��j�|�{�*۽�O5Q�`�ۧʲǙ��P\��"#�x�^�()l�̈�i_W<
�Y9 M�K �,,L~D�{�&Z�h\6����σfd�ha�\���W~o��
t]m�{��3���s��}�ƣϞǴ����F����}O0��y��s��U�3՞��(���~��|�[乍�U�%F�d�vO�6B~���)ț��ů���G=>�r���>�����=w��YN`�"=E:-,����{5��q+��f�<G6�c��9��w�P�9�++���X4rS�R��Q(jOjWk���Ý)��&ܯ�6�=k�7�c�"@T�m���wZMt��5���Q�2d��L�9f��0�����	�[:,e��"�|bS�n�����ś_}�S����c��o��c:k`�9�VQr9����X1-*��C*�Q�f�j0����Ҽk"�yL�ݐ�Z�g�c�^&�G��Jl�� S�R�u���T}Cr|ŵ�|�*�w�����D���8z��Flf���ƣ�9�S>P���f���L���d��`$�MpJ� -�`v�,��X��̉,�����g���
nF�=~�0�?��:8����=��
KB�� ���9�6�\7%�6���Y"��Ú</�*`�
�WrD-$x4�e�|h8F���=]+�\��suʣ5W���'�{���)`A���:�$����z��	���_��SB֑�Q���en�4��s<�ZU��1�@%�b���>�`\s��Vxp��g�=O`�/�&8!5fXq=�Jz pk�g�����9X`o�ZWUϹ;�*&iơɐx�7�&Sl�:��ͼ���U���)�N.�.����z}LX1e�s:G]��V1e�'���1�X�bZ� `:Ĕ�.��qЮ��k����-]��M��Т��{Cɩ�� ט�R~]��.Yfp�5s�Qe��5cd�z=��9fb$�W��+��&��X�`?)�r�[
����ݤO���Z���90F��h�������9^5�K�g����UTx�Ⴝ��� z�0V(0Z?T�JοF���8���$�VVH�3p$}sv>�)���U���яF�H��������&	$q.+��M�&�؛�����x�]7j5e�&�5+V�]6���_>����?��N���P�;h�;h�Y٣��RF%f<�j�h�P�9/�����䊣0���S�v��Y!54�ck"%)K�CU���HJ�`ZR3�`|�Q�0�A����<`���r���p�MW�G�z^��[p��&��M���ڳL�<1����n��3���tj�G��>�z�%�x�<N<
/������cV\r,��u�� ��٣�h��l�����F��~f�T�������qNR���cg�W���-��HZ[kE�,�BFTh?F#�=ײd�������Aa���S��w�8�Jի�#�y�h00��� ���I�~�eJ�9'	`g��K�u2u���!\w�1�t��xō�RE��C^Va=)#⼋��B�b��x��~�	|��'���_��}̫tE�`��FKS�v��Y�*����Z��������E�*�@��CoW��0�s����ޟ]�����f���(_��RS62�����E��}��Glk��d1ْ����p#��Ͽ��eM�K!짹%%����ן�����ό0Zt0�V4F���2`�Y�|+�⎗�}奇��Ox�(���p�sqs���J���wn�a����^���nl���o9�����#�O����x���=h�c�Ƣp�cTR����_�,1��8(�l���c%T�j��K`��h�2�b��yS�@��i���h�x���+�-��j��3T�3����0��0�NQ�D���f���G�?Q+� 0m�sTn����6<+"ϩ,A#��k^�h3]��ŀ��ׇ��L��#o�I�t��c���x?�|ۑ��9�V1��O>��|��8=kZ�T@'����D�2�P�-�u�mj�q��c��W�^�}�����o��K0�I��xjbl�L���r��j�sӃ��P�dO�T�w9/M�w|�U�i�TQ}L�X����o�d��{��X�"N�GN4�4C�Ks\Zō�����˥��KY�j)OU��-�9����J�T��+�;K��>�u����H>�2t����ҏ_��6�[`Q��C�@*�1�f�#�9/��荈�oW\$���/{q�H�M%(]Y]U���J]*���	q4��h��q��z4��9���a�Oê�8&db�}M�(9�-�	~���3�1b7%�b��
�&��Q��[[�5�p`�K2� .ñ W L��1�v_�Q�K/U�����-h$�U뭇�ݾB_���k� �s�s�W2��c�3Ȫh�Yu`�=r���;�q��t��Sg1�E4�]t�}9�)�da.6�w�b.�$����r���O'sԘ�s\�JK�&�S�8d��S6����p� Α1$"q�+��y�Ҭ@�&�/�z<�$�L�?x@`J���r��S�����"�_��>[s�����!�\��4TQ�O�ݚ�D�֒�iJ��ƒw9n;��V~`��������L�k��"V�{0b� �Z E1���E,�>�D�r�ks    IDAT�4%�P��o�.��J	E[ �'7�aʁ<��8i3�
De���39�{��ZV1%gl�O���Ho��h����So=~�]o��sd̵Gb�Q���o_��|�~<��ETZ�P�<�,G��DN�G�|
��I�R4��}xc��=�C��QGL(IƆR¾���f�s��S����Eh��`gw���Fj���5l��[T�_�^�h~�|6��k6��bL�gO��+����2�z�u�����[�a��ߌv#�
M�6�^�&l�ą���N���/���'^ƃ�~O?�"Ξ��dB������Q�H.�5�1�[�SL�H�J��K��������2(3��!��35��{G��<���R6������ޓu;�"�m�c�x+�O�|yN���m>5�����)z�:��1���r2Ƅ~�a-E|0��l����^q7�p%���0���.;���bu�ʰ����,�Ƿ^���U��;:�w�ǟ9���1<��x�%��0�6	������9�D��K��8$��z�,��ʉNZhNXT�l�yv�d�ޏ��w��t�W�L�T��Ho�Qv�0H�]�#{�FP�d�<� �&f��d�&G��þ�k�~�G�ć~�Gp��M Z��
���Ii����<�?�����)����**��26)����rl+��^q%�U�K�bک���#<L
ըR�<���u�V���b�B>�9�I����6"�*;�D!MU��'�1�;Q*�Kg:�ލX�اI!6:�S�$��41��-��N��s�o��UL��q�Ӟy��D��H4?jx���WQ�X�q1��<����J��j#ۻG��f.��DNOh7	L��:wí��y�4�t^���x3���1��8�=t��9�J��M�Q�ԭI�����\yY1��O=�?����종�WL5d�ه �lB��C�����:ʮ��bG��?��Y� +@Կ�`���+�z�^R�N�A+����M�O��SF<}�s�]�d`��X�X) Ϲ��_�c$e�DL�&j��nP~n$�%��)��oZ��)n?˗8�gh�Z2�����LSγ��5�W��}L�%������516N@���J�:ރ3nQ�Ʋq<��Y�K����XnQ��to"��A�}��F��QV���*1�� ��Ge���J_��0��Gl�I��着���便������.�Ԇ�$�&j=*��iP�8&s4��%Lo�����τ ��g�;9�2a�,9��!S��E`=,I~�t���`Y�<�
[R�B��_�!�c�/��� I�QȽL��D�tI�m[�v��z�f�>��]�G)�%0�9}㝞�Iku���Qi71������ӕ��b����|��Q��t�����
�n~DVQ��s�y�bD�j��P?O`� 0�29�9Ͳ{lH�QW���@���s�4��&�0��I�kbLɫ�Z��4{jէ��"��'�=�Veb�'(�1]:���>U�jH�M~d�Utk�:�I��L]����v��X���A��$)i�(�l,�ź�x^,M��q�&Ф*}ѻ�W����e���r�hĪ�ab�=aA��4)�H+Q��L/����8ݳ�Vv��ps0��{5���1���!��!����Gx�=���}��N��qG]ig<����G��y�Y�:49��<�SxQE���
�DB�4W�4�+@�|�2����Vы
F�U���Bpgq��3ɻW�\�e�;�p����� �/o	D�}L�n��3�h8��JƑ�����	�;��x��q�����5p"L��G5�G�����e4V1��@��T���K��q�������O��Ͽ���;�ޙ`��Ɩ���2�	d�R`*�}��o�wl}���U�ZE=Ē��TIa�-F|FT�����A�^<;��!1�C�z�|>��G�rг��j�G���3�?|`ꓛͤ��{XR���ڜ?�?#VT�h42�ݷ�ˎ��7^��n��\uW_qG��m I�%����W�I	�;�1�6K�[3`ck�ϟ�C�<��=��{�<��tB��}�3�����sM&��H&�TZy�'`o��$ٶ�h��N�:In�g:i�KW6҉�����+��-w�g�Z�<�E>&�+��*�I�]�ve+�cNu���:��.��?�6������=F���:a�As�}௿�$~�?���$QW���5���7�[����eik���1�B��Yy'#v:���rK���L�Z�$w(���n�9��$l5ҽ���@�S�Ic�������qnj�,��8'��1�~�)��c7#��|���� ɪȺUL��{(zH�W*XiY�t9�`��y�{Zs���h������H�<B���Ou�J�zT9���%� ��c�:���WR^j���On�D�L�&G4_��%�n��/�Z�]�Z<��3n�'�0�e�֊�,�f~T���?�����h�0`:r`���z��_��E�]y͉�L5wLsK���n�Q9��'~>�{ˌy�b�L$�E�-�o��ސ�-Ŵ��n�t�U9��[��Y�`8��M�=��Ѭ�*�ޫ�`�e�x�MتMv��6�y�b�̴?��q��̒��t0�&cF2�t$���Li~`��5P^:N��&0����$nF��(Kz|�KO O��m�d"�q�0� ����d�� ��?��X(Q�I�`D�J����Vb�q�@�����B�Z�^sߔ;[��z�P�{6���̭Jm�%�ub��f]���q;ܴ>lܓ����~ό�L��Ge�Ph_�iV�0Y{�C�h��8��C��[ mv�Z%ٴ���N����s�<��*m,ͥ��x�vx���ޢ�H�uȹ\2XvW��G�RPg^�.�3����H]�4�LU��Q9�I;8s��d2E��E�ؼ"`R^�̹!X�iU`[,l\�N_�rNp�}Aq�*��ǐ80w6��0���j�q1Li~��i�Y�n��d/F0(Kv@��P�&��w��LSC��(b�yM4Zjfn ��Y%>�Z�=j�,A-�ww���}�$����<X��*�B�Nl�a��2^�x�qr5�x i��\��A	�F��-��K�i�S�9i��tU�� �&D���i8\ ��	����q�@�"v%B��tŨ����-'�"Y5�����2����z��c��8�	��1*�����Z���W�U���T���p<{
��?�>��G0��Q�J��R�Fnrsg�#�J������S�����HP�)�pcH bt�J�]���R;O*��]W��Jj��D�
�Z�'��q�*�J�IR���
�.5_��Ͱ�[Ǎ���\��:�#��p���u�ܶd/�TT��6���1[���>�[॓;x��'�?�Sg�q���7F����QL�:� T�k�'/	$��Z��=G#����Lk�B�Ǩ��L�Z�$b@������J�X���nڈY�o�ȱ�2�I:vҽ�`U#68����C�t*��	F��X�{�ay�T��j���k\u�e���+p�W��ġ�t��.���>%"A���c�y6�6f8yv�>����G���Oc{8�t��"�K�K3�'I2�T	xZL7Tf^�W�"��S~dN[?!����),�D�)���F`�'ì)v�|�m���~~Z.eU�Dw�ZS<v7���E�[�L�q��k���}���W�@�g�ZM1��s;�'�~�O?�ӛs�k�/�h�W���{���nY��g�w.��\6��~eT}u�<u�oģ�z�=c.�-�0�,���wĈ6�}�/�v��|c>���
����#������8��k� �mw��A�#�l�x�k�:MS���rp4��zLW�M,ULǽ�*��G�󌅙|70U��|������h��ƽ�`��	{L���a�mW��>S��b{	0�����m�h�b����+�w&������̆+���|\Le��#�)��o}w��*��<��5(ΐJ ����w�����\y{���8�6P��m��U��-NL{0��ؕW�+Jlф\/>�`U�[��������ԆW��8rpo��6\u� Z�EĠ\Yb�Y@�}|�[�ŉ�a!�pʓ�r��F�]U�o�|�<�>Ɔ���uZ��H���6��������h��L���L��ธj��*��&4�`��*��p^kM�R'��:,�	kac_:��g�&���\<��v*Z,�.`��_�-7��g.)`ĲR��;��G��j�`�Ai[��|f���Rv53�m232�5�'���9��ΌS�+���%����NUFI��r���y�@S�x^KrY�V.�.��U'<��E�T��0����1?�c�xV�r�M��$�q�������s�zu�ֆ�6Nɞ��`]#m����f5�b}�������5��0���+�p�I`�j��s��Q��h���u�@K9l���w2��x�;��9ri���ΞUT:-T��4g@�\T��9_�T���3u)/u{�*ظ#��4:��]J��YZ!�-U�x-���|��FG�%�$i8��f
���$	��,�o9���t�)f��J�Y�1	���)�3&U[Ix��5�|�|^J�<Q��צI�/��G��[QA�=f��K�	��J^T�f�-��O���A�ud�N�����#��n��o�vt�����2;$C�j�����~�Ce�L������i<<S,�[h�wp��G��{'^s�!��<d�ʢH� t�=q���z�;8�1C5_E-k�u�f<t@�$7�FO���Y�0-��0�*����0��J�'�J2�LO���*�j���J�\v�j�J��!T��gQ�R�9d����u�댝8E��V[`>hX{�c�[G������ǭ�\-W�;n����p-*C$���ʹT`�]�*u"lL)�vt����%���Y���y|��S8u�<�_Xǅ�Ml�͖��"�3�RQ��Ӱ?���|L:��X0���zQe$Sl[�,	j�WS�F�x�;}�O�f)�-&��[��Mǘ�87����zCY����E������ὸ��!;zG/ۏ+�Ƒ#�q��V:4N:ć�*��~(,K,̠i�� ܕ{��/��G��SϽ�'N����1Zd&ӭ5������-M�d��~G��φ��>�Z�����u�w�+e:�HD�Qz����
G!��#���a����y>c�Α#>��Y��-e����,�������7��q�Y��x��gߎ���&^E���[BG����?��7�����7���XV�����D��{��L5�����m�>��*��T���J^"a��I����E��
	�d�#5A{�{KF�u�c��(��$�7�};\�,�_�ag����T,��E\�\�{uag,��*ﶰP��q ۢ��&����5Gt��t��38�A��|m�������"���9�j�a�t4���������.���ò��D�k�dY���8V(����6Μ�h���/��^��R�d�5SmjƱ�[��Ĝ����⸘l1��+���7?��o9�9�?������������!�U�"�0�U1-$��Q��d��r��]kɀ�H <�H@�ج`i{>���(,ڍS�ӬMq��q�=�E#[bk��<��ֲykO=w�x�	\ܚ������ԁK)o�XT����+�����'.|�2��kȡ�
�Lf���$(B��YS&.��4��5�M��:��)�\�DTm����}IU�Ê��Tp�aɘ/{���	P}��=!�����.��q3��I��gf������ؼ̒f[�Cg�.%�L���^A��N�G:�M��Z�ZNb�����F9)��!���Q�K�xm1����:�
��K��!�^���k���N�v9I�B��4<�~R�x����"���>���[��~`Fe5�d��Erp>Uo�gSli�t�7�H���-Y�5d��f�>%��3�VZ�P��a��-@�`P�kL&�>síU�{ְr�<J���L-��
s啔wS��=���V׺��RK�>�4w�׹H��2@on�6��o��j+���/����{�~x)�"��v��o��2��To��b&#"i	`L9"��K�Q�'`�#IŵD��Br������9�f��ei!T�!���}\D��L�W�PY) w����q�(����Z���^ĝ����ZuȔ�K0}�)b��.���wS���|@\�
�L�iKEOR9y2�r�w�шW��
�1�rn:��݁�GA�ٹ�j��b�ٸ�h���[�؏_��O��2��T��q�����O?���c_���i�"�ݽ��sK��G1]O�$�M�wahO_w������J��]�흛Z�������V�?)I�#P�Y��܇ʊG�M�o�^r�w�2X~���$�t�:1KY3��U��,&�v0�oI�H����&���2��=w��;o�G�hӯ#��w�nMղrb�S�w>j3���裷ӟcs����;�6�z8u�"��,^x�N�Y�鳛�y�4�sk��	�9n�u�x�<ڞ�������K��& e�,*��|��=y�z0<��/(�f%T#X=��ݪ��ɰw���{W�w��=+-��k�:*Pz��~�����[�BZT���'E��L�g�<k3�"�r&����G����}�=�<���9gQ�'!�<[2ƛ�+�tUV�NF�D�vkc���e3h=c��k�Xڕ#��n�+-��o"F�괜,Z�J�ň�47yw\L`9I@�g� ��"�H�ꔞ�$娰���}������G�?�x��V���<��O���FG��7�'�U���0�v1Yҝ�#0O�D�����p��:���|V�B�C�|I�N!�@nr���d^8���d��]�97��LÏi�����A���<�
���Q�k-��5p��&�-�G�s�W�=�h;+�}nX�J*�2'!����Ia�j橫�� �r���p���gA`*_�
L뫫��q1޾E2�Ƶf�}�N�Ý=���+����M�ㅔת�y��n���z=���v_Ĭ���&�5`VsrG�����i�n�2��&"v�b9	�VG�8�e��C�������ӱKy����}�oq+�W��q�u�S�G��h�irhv��ǥ��lI��Q�(���Ub�DeA�H�G�,E���0l!��Ш�p���*Sڿ��2Go{ΞA-�`��5\}��X;p�Y?z�i������R�4�N!�+|!��缬���f��bv��x_�:�o$OeFZL�^Ա̹��4��&P;�b�bI��%@�(I@�4)�����w�3�F4�"6���kRc�̬�֕"]h:h��R<_��%c$�@�=&尃��~�X:����`e�SV �mm�`8����,����`��i�Z�k��di*Մ .�tL�ыJ�X�#eu��nf�mU�1����jy�=au�K���t0�ˌ���]I\0��|�P!�-zv����Y���M�y�=y�^Y��-f cA��b�岜גND`
S�1���@+%d!�� ��?�r�3�cg��=j.s��6z5���D}	�|��*���D�"]yk��&/Q�j8�Z<���z]W3��0��/�nst���[J <7�C{Z��Z���FP��}�d^2H�]YEA��o�'�笫49)f5�7��%5����代�����t�uɺ�/V\�}PO:��Ҝ����H"1V����ƹ���Hձ0��KM��m%IΥ��iH۬�����o�k���L5<�r��r�	������K��:LK[��nF�:��ɤ�����{���`K{2*�Z�>��s�*K9bNz��h-���sx�ݷ`_�d�̧4=��s���lM�/|s���ϟ�`�����&LDI�գ2dU	]���gs�.�I������s�:v=F���=���F����HZV-\��q��Kd�b,���Ҍf� '���b�>'�jnu�A�)���Dᔤ��Tf���z�C�Z������7��~��8zpM��~��o���0k%a    IDAT���W�~\���e�Q��G@�P���g�G�¹�[��q��m���7�\%!5�ً�>?*k4W0�~�W<D����ƒI���cڀ�l�f#"xvQ6��WѤ�f3��V]b�Z����������8x`M�tm�ƶ�8#%��{�ܸo�޿PD,4� �z�"�M2}�B�>
_��C��c�����iMŃٲ�"Z5`�5,o���>�*�n �����.���4'��4���}6lIyR��\��	"W<U���3�
���T)��+�oU��*J�9b��U�ޕ���ڜs�N�e�
)$&4S�c1�B�:�[�����+�ibOp��ut��8�%��9��_��?�5����ek�V�3��nʳ:����(��&֙#���jUs`ju��GН-�����"���|����4��1�H���Gh�i:@�ͩ��j����oi���@�?�"g�=���	�=G��Ĝ��
�t�O��8)͘ L�Х��N�,qp�},#?�Ǌi[���@�C�}�}�3�S���Tm4���O��q�K�頱�zL'r�-��s��F=UL�/\�`��t��*���R��� ���L굪�Z�Y��ӑ�z���J�fÁ)+�<g�ى�v����-_�R_L����q�;ǿ��7�W�T����2?�#�}����_¹e=�$K1`j)�69M��By��v$r����rI�"�Z�7 �j�Y�k�y�v��9���c:�Ĥw���~����[o��9��	��?�/>�E��}��j���ux�]oD���ǟ~O�8�ɢ�e��	+�D'��ʫ/A�U$Ln=�{P�����E�8;�-Ȕn�[��a�)_��>����kVIjXNZ�����$=|���BsC�F`�7�V$�v5e9��q���|ݻ������/޿`��bN���Q���ȖT;���B	/��d6���6X5`(�P���l����f�SJGJ��ٺ�$��J���Z���*�6��n-N���/k�}��Ҕ�2������H�?@��%�n�d��𒹈�pa�j�vMJ�]� ���v�w� =h��"%/�x�k2&�wZ~h��.�u�׺X�8.ƌ�Mjd}:��hl�h���g1���}��ۇ�#G0#H�Ym�D������f��X��㵔��g�#A)��ɂ�Z��4��ty�K6/�f�.�UM]�c��V����֋��h���?דn�ͪO��y�&;sߥ�����:�.p��U $��9�)T�l]��1OPa�����F�V�s�����b�Q�]�0j.1�S��d�&�*z�c^e��&۴��0���#�J��,�܊�2-{֮����Z:[R��![�-���ÿ�
��R#��a5��R��W@i���ʹ8zl-��5.���)��H���?O��,�=,��8ح��}+~�ͯƱ�fXA0��g��(�s_;��|��ƣ/c�h������� �W�2��@��pg	��+��Ǟ8{R�3���ra��N;�޸�'���,Ϥ��֓�q"9��OF��#;^�v?��ɱ�\�P�]5R6��xńj��{���E�4�f:�B�>�M���n����*�t����}V��Y?ί�k�3E����+��sWfΧ��We�?X`<�YR<c4�h��h<��#9h��&�|��h�Ʊw����\���3o��V��o�TԪ�8��dh�r��Z�Y�v��kU ��̰ڭbu��ߗxo�1��X��d���m�ٻ��g�?��x�<��{�,.n�0����D��&0Z�5�W �:�*)�:�~N��JW��m�#�c�;��'ͣ� ��83�8:��r�k=���8��n��-���f+h�����Z�R��ubF����e��喺>����>��g��`1^��r�Ľ��g�s7�<\A��Q�b��ϫ�/�����"����5b{	��;��-�J��q�O����6r���чf�d�@�($ۡ��|tctB�L����y��ɔ��H2u�@xߧȪ3����G�oWq`O�\uG��e������X�iJ;ݐ��i:�a0c�����-�9���Ooh��8�hA��FZ� �H����Y����s�X0��i�d���1�*6��e$5�NH��D�*��-��6ΞǄ��TJ�����Ƕ���TO�
0����j�)�����C�E0ݿ�N��B�MUl�2ϢUW��4ǔ�
G�q�í�n�>;V�ܕ*��pe�O �[��;��������qS�)�b+���~䳏�w��8�hcT�bʚ���-� �d{c��-�`z\c/�؀�%���@�'��������A��?Ǝ�0\��s�Ư��x�5��y�pq��������??�!#�hvx���=o�=j���S'1����9����UVWu,�m.��)c,8�d�.z�75��H�RC�kE��ꖔ-qƥ'�6���
u�	8�H���?jI�[�Ge��o��ƿ��`��9*f����d��"���OdC
�ew^o"��]�+&��@Y���r�`]�-�́�Kk�#V�(M��4&�����<�	칆��QZw��$+��`�R������E5A�5����c�#T���;C�,�GN��u;�dl�`���:�o�4��XE�7�m�Xň�I�OH�G8_�\uKϬ,c��(-�'���&�`l�:Ur��qUKb�,����
��=�yQʊ�'�)%�|���/�0%��f���Q�)yU��F�șZ�%>ӠDxkG���Cڟs�t�g�N�*��,�Č-�~	�VxaC�LY1`�(�A7�Js�c��Z.K�DHg$�$��7�$��b���@�
�%����$_1b#d,��N�������XNfr�e��L�o�����$ݭѫg�櫵M��� ϿVH}=�J0���c<�z�ԓ�U�0��8P�f鵕��:�d'�`��Ƃ�
yq̢K":�m�l��D�i�dR���JO���^߫�R�t@����m=����V����BNi�4bOJ�4�m6�lp���������O�G���U����s-;3��OO�����c��Z���ّ+,נ\^�k�g���bF���$Ӫ5��������)&�\�F���B+W����Wp
S���Lب2��`�����&?A*�GI��u~x�_>+�����C�"��S]5�l�� �q��&���us\}� ���[q�+���7\����2_�U#�JU)���2��>i���_���`ˀ�9�d��O��*���B���[mi�d*cOVclM#H��<��g-M&��#����Ŵ��*އ��F�z���B�L�����;�9�����7���3��'��S����h8���\A-�r����&(��i�J���Z�K�ECc-?�f4�î*r�x)榑l�&3��X��H���L��9h��K�Z���l�e5卝��g� }�gب�ȡ���T?�X| ���Q��&Z�1n�j~���=�9�U-�e?�m����P�������#ϣ?����U�@����)��#�+iog�=�C)1<�H�x.>��@W��x��m����g`L����j���1�������=����v�r��8��݊�l���K֬��4B�O�����䳧��/=�Ǟ=����eS�f;Qs܌,��v�&��!�՞�0�ET+�ph���}���6׸��`���2?�d��J�^�1�4rfR��@s�jU����? LقɊ���uژb�����<[����j���.�9�ـ��X�[�T#�*�p5in����5�����l��c�4[Q������Kx��{U-��]9���2q)�G?�=|�Ͽ������VL�q̥PH.k��|�� �����.C9���%�5��W?��"�B��j��Y/��>�n|���:�sQT����?�Y���op��y�,V�n{������2���3x��S�;X�=;4u�A�z܄�+�4&���.�c%"*�e���n�C<�Y%%K}��-)�1	����er��<�g�r�GkS�c�U�����w�OP?0��K	STz����|/w�]IAi��N(�'.�W�'�$-1�z��8�H�����u�V��X�M��w�ͦ�Ki���CT9��� ���r^�R:�yk僀�c���d�Q�Q������[����><�d��4wh���ۋK��;b���FO�$�����^���z���ʷ���yW�}�k\ � J�˫9v��*]$���6�e�8\#�R�4��Li�_�}�K2�3�d�5�d:��˧���V_Ug�^��Ӭ&�fQ�90%	d�8�(��	Ҷw0���l4�����"iK�b��ꬫ*�${9.�⦀)�~^�HV�\jL�+|�I(* ��+N����$Q���?Խ�a� n`�`�9���G4XJ\,��X��2�&���S�g�u�'2a������:Ib��w~�GS84�>�բ�@�)2�coj����1#.	����ׄ�z.�Ծ(�3I� 2�ת���Ju�Y��2�Y�cs��햘�O����֦ң?�w;�� �g�̱:B"�b�$��Q�.T��U�[�6Щp�W�_��/���&_�j�9��l��/�g_��>�u���Va��\�5TTdFag��[��T5��g���*�ך1��kK���Հ�zLݍ9�{��j�(��?I�$�����п#.FR����L%�ߙD�Ia i��M~���n����z[��0�����63��_�x�+o���_�ˏ�ޕ̪�U��I�*U�=J�&
r'�h	�
 �����<����8M���=����b�v	!��/��X^�N7�oJ��%yj#���8z��}���ȋC��
�x�o/���x������'�����������+-���xᤄj�i��,0����ƅ��(	K��i�&���\*D+Ai�\Y�o�5x}N�P�\aО^䭱��lΞQ�(jF8.s�k�Ǥ��	M#�����G�9Ȗ�����Ñ�4 n�ƞ�oz���{7^}�^���m��^��ϟ��π/=�2~����C���{Q�9��&�'��*M f��k1��)�s�s���{(�"�����R~o��ʾ|F��p�Y��Ke�Ze��Ɇ��W�wߎW�t�˵W㸳|7y[����h�.~?;�����K������ę�9v(+�L9jF�.]�6�0��n�Lof��Z��?J�i~����(�e�
uPCR�::y��2/I�;�ͥ�����)����AʵWUL�*���mM�`AcuM�G�n��L��ܝ��꫟ϭb:z�vdŜ<Gs����Mͫf0�T�m�R�pKM�`S�����O6���/����bZ���`�J��x��c�Ù%+�+�/L�K`*YVH�t�r��Pc�+�(=���d��,�Ic�����+z��U�h�����7�o��O㎛�I��0�İRŷ������x��G-I�.p�[�ś��.��s�>���=�"f�5�%Qf?��uڈ<He���XZ��ķ���[;Qb�j�DK\Y��3��^n:VM�L	xu
��̬�u_��������ד�hQ���F���b-�W�B �a0t��DX>#�`X��*n{��t�I\��^�Qi(̮�G�&54�-�P�ԙU���\'��'���Gs"J����#B�j{B�[$��>�p]���2	U�_{7���-:����nn��DL9�@���Y��Pnv���F��X�KnU�4Xڞ�ٙ�L�J%�q|ʀAal�%�%c(�� �$q@_T����\ɪ��t����:��(U��}�����;���o�g��t����Q1'ZŴI��V�����=]�>.fVeϫɝEj�LML��tta��@ @}������A87G���)h�`fi��ġ#+��|�zY���0�7��}��b���x��F�V_�,:VJm�-���/����3D�qG�H�8t�̂�H��&E5���W�S|HRv�� �:�t�ɡ�S�k7`��-�a��4����%w�N���C�)�ɞ؏��Q�{J���8�~��\Ҽg��/Iu�����5]֥sQ�"lw!����yU����4��Fp:`1�D}��7��
���~�]$����J�N�����_�<{#�Qk��P���RM[�>Ks������fU�ݬ��"��p����Jga85�Yo�C~�xE-�Y�x9pKd�ߥH�w�����Ϙԃ�}뮺�*�]��N�,n�zf���y��i&*���Q�� �!}+���YL��i���8~���\~��<{��!>�bsSc��#O�9�������`+��%rZ���-�f�y�;A�V�q�t�r��,N�y5����E���R�c�D$�WrF���c�=w���������^��s/���'^©�[�v#C��@�ݕ�N��j?����G7݆>������y�z�ޫ�k��rR���WI�S�e�p�oWw0��kk_���~�p�wI�%�oi���
�*W�.�f��ſ�����H�|H��0^���u��w�����l7�p���^N������9<{r��~UI�U��2>�q[�2	�bDb�aX^��z"q�v��
Lǋ)ռl��� U�*gBJI&eU<�Q[�m���k����Z�����.��Ȥ���"�ݽ�v�R�g����	��G6��ă�=��QUnЋJC-DQ�R,��AS�""���J9K()o�.O�Jn���TS-�丘F^�몜r2�S�;,��R�X��H��5�.�k�����6�É�Ѭ��{L�MUL���J��"n��q3�j��@�t<0`�z�Ξ5d��_�Ǵ\1ՙ�b��B
�<J�G�/G�W�-�~�Cx�uk?\�ˊ)��`:oa��`F���+*��j��i�lE"!B�gv��o�6��S-R�QQ��j%�t�fe���)��Λ���gp��$,��:��pz}������矼�e�_}�z�=�����ǉ�O�;�<�鬍J��	�݂ �ɿ1q�n���?�3>hg�o$v,�`�Kɡ�[l,�����f}D3�����3IzM��>�N�1��7�SUr�J]Z���D���)Bg�39]�]jQe��Sl��E�U��E -�i�vFOm�WA}YV� �U�>׀�&u�ͦ*������i�|q�ǻ7�0��5�E�<��|��.�go��	��8�DXH��g���oAX���ں6�ʇ�9�01�p���V%R������Y�o%W���#K;�{�+���~���Lwɜ���ޜ��[ۀi�Z���,W��*�g�����'�t>&��&�=e�4��ڳkG�a�gV1��`n1���i>�a�纾��)�O����=r�^b�\HGKa�����_����QKd���P�k��}uB׮�����1��'	&n�F]s�dh�޴��6K��I3�@�-0:��Wr^*F�J��I����"^J�2�Xj���K
E��G))-)<l=��*��0
�0���y����-Mq�[�|[T�̈U+��L��e��8���S����S��	��$g�Gk��+����U�8������a��J�?�៙��d&�|yS��19#�����6��n�r?��{ބw��J�����Z�D�9��x��1>���q�מ�z?�p���
j����2V�l��\�%�{:g[�Ɨ��E�S�M�s*zZ2bq0E�� �K'B"(�K'`�S-�8ʅ41^�{� ��+bNfv�`ο���cD�޻��V��i�'�=��S�A3�|�{����h�D3���5zO`z��G�[���/hݷo����Jm�湬�,����QU3���_Q��7k��{��QL���7�H�K>�f���T��\�����e�ƽA���C����1vzc�o�������?�g�}g�o�7��s��c^͑�VPkv�������@�����8!)i���<� �hĄ��U�]��M��(��~քI�����^~>��cS��Tϛ��0s��{�?<�^�Z�.+���%\���S{F�@�    IDAT\6B�W{�gsPΗ��t�崏�l7^�ů��=x�=7b?�^TI�k�1T����@�}�����N_���؃��~��֛-��Oi��vI�b9��R%�P*y <�a��9���DYG�Q�#?hy�M~Ζ�_s�����֪x�����o}-�������/������ދ'��s�г�����灿����|�{5L�ƈ��v�%�Ai�򞙂JQ��oaN���$	��UJ0�����]f͘Ԩ����N�SL���V��Q S���?�L�♛�T������ƃ����Ǵ%?��״F��TL��y�bJ`JϐZ����U��T��x�R`jd�IG�I�d�|��i>�0�w��A����A`��̏~�q�����y�J۬�%�r祐�F�Ё��T��W]��K��7��_2���nleB��z���ᶐ�����{��?�G���W��0�a s8{z��������t�^~9&���=s�E<�س�M��7V0�A͒�f�l��s1c��.4s��8
P���PdY#d�z�{��RF]��C�U1afo����&k�����s,�k�U$w`�J�n{�GŖ*�8 u�ت1Y�Q0�~��хCg"����*Q��ZH
-Ep¯��]����<%2�h�Y����[h�i,Dkx3�
c�s3KIݯ��>�ٙ�ְ/Ìt���팧��T�4Sg���H9I^�в;'7ik�ϟ ��R�m���f@�$ۃ�I����%@Pp��^����t��T���'�Q�d���H�}ATD��%��tg5;�cE�=$V�o�iI�n�^�u�ڠ�W=[�	6^:���Mp�Rg�>t��Ȁ)���Y(��e����N.n`:0������Q5� �"��*��"�i4���� �lϸ�gJ��20�M������n��0�� ��$NZL1�T�*��~�~u��{1f7����Jy���q0e��B .{ %@ڿq�D�����%�dT�=��@	i�ׂT
b*��b�k>�"��i�g%�$�E��2A ��
`L}�GdY�Ć{G��.%��KF]^�H*��t��;�WE�u�_ŉ՘��{����cz�Ŗg�2]e{A�d\D��9X.�`�S��0������w�}?���|�bu�vU��\����i�������1�5Pk� ��f�V�̔ثŘ���TK&~nZa�� ��vX��jm�ɰ��Ɣ�1b�6���oe�����lΗ�Q�{�RI2��-~�I�`�<�r�C�7�2���9�Ǫ�bē����gm0@�60�m`6���?4
�k�u�s=r G���W_��o�7�p-�oQ@"'۠�t\�H��X�e>���FEu�)�␈�	嗎���7Ň�W�Lb�p�w���x�x��p��y�[�w��<�s��1����@-��BY��m�V`�0�Cƀ���h�O�I�U�,��=�j9ZM�`��0���WxV���A?(������"n�M&��3������q��;��wň v��MQ�8��֢ a�p� ��͆����9��0l ��x��oį~�ݸ�#"�(�4~F��mI�w��SS|�/>�O=�0�l.�OZ�W��tUɶ1)vM��<7�8��Ђ��c߇i�ٳ(��D9a����5*ܔ���4YՎc�1�w�����3o�[��h�[�f��n�'�G\�_-�Iz����� ����|�$�۟��~q�eyg?FSz)�\j�`���<0�v"7�"0���=uVY�D�z��2�v���� �6T1�Nf���i���^�.�m4_R��@)�J=�J��2��wa��-Szp�i��>Tۭ��HR^{&y���f�zL���=�Q$%i�^����"�9.F�ZovΨ�S�5N�nm]R	�������g�k�YS*����Y�}�s��?����)yU�/����X��T�L"�Fr�Β[�Yp��.Lr�3ԤA������i��d��x�y��9�m�y�����gq����٘C��)pa�淟�7zg/l)�t�+��|��O���ulo�P��4WL��ڔ>̚��t��T���I7;p΀J���@��(S�BFV���xUb������,v#Wb͆b�l3�Љ��t�l<C�C��_����|#*�.*���%F�Tu0�+y:�-0���NHmC�?0v!��$%�E/���iS����aɴ���&%�(y�j��l�l\L�+�1Ae/��a��pا������g��mm���{��W�}ۜNZ�Ӽ��m��iK��6��R�	��e=W��[�D�T�$������i�yTk�	~��\H��'o^�6�H蜵q �R^?�A�E�{%}�,.�5}��t�.�~��)e�tk�E�Ƚ�{Ta��d��;c����^��^Z9p ��.Äm��T4g6 ��r�4QE>�a��c��XR��ꪀ)��8[K}q6�� �Uj��� J`za�^���s�I>�r}oF�x�}H�pv�v���<C��l�L�!eL�ߟg�2���ܤ�S�3�	&�����K�%wi<���"<�]�TН��/OL�ɳXq�uPUS��#�>)ъ=�������"H�����C9>Z<
���-V�RR��+��<���R���b�o��|\Ȧw�KK�.A�rb��*�2�%��Ϯ"��-�uc��Sʉt��.�A>������6�w��@6�ď��x�O��]����,f�����k�cώ�_?�W��7�B����zG�����f�	�eK�55�v��ԝsF�HJ��3G�3j'I`��n�ʥ�+�=��o'!2[5|��Y֖a	�Qe.����+2�'���9>�G������w$p�M��Y]q��{��M3R�1l�`�2�HM45�}�<~�/��\y9�>���+h���A��Z9%�4/b��ɟŃr��`��!��cJ�����xP��Y8�db;���t.'`V��r?�.0��������|��i<��	��1����T%ju����O9ӄE)8έ�F�^�![�Xe��&�ϕ?բǙF�\_$}i~��dJ:S���<��u�U*����}�Y��ӹ�?�~I�CŖ�?�5� vǝ"_�k;��Nx�)eO�sU��\#hM.���-2ﳜ��hܵ�����ď��j��~�]���Α�$(U�Y�ޑ������/�7�,X���f[D���RHxb�U��a�`�uB"��ww��.!�
"�XBS�ZX�w��H�U���`Ux��p~����e�X�E,Kv�/������������	���sa4��q�}�~<��l��\��`�Č.u�e��z;c�HeG�*��)��2�Qgi��6��:f�	&2{�zL�VPir
�b�d��:��v�W�u�f3�1�°7�bQ�9��	L�����>6Qp��Z�-Jy�����8{��H9�����b���*�ɉifI�z�T�ȸQ��{af�t����,����/��kV80���=���pz�BM,9C*�'�$��&��h�B�d�Px�|8��^��-U�&�&�.��h�"05��L#�'m�>:+u�v�M��'���:Ԫ9.\��3Ϟ��� ^:uA����Z����O�ث@���d�rwys+;�X�]Tg��|�hu��d��n�W�l�Uŋ��:L<�J>�@,\��q��X����1]�A7����Y�-{L�3�yo��,���m�_c;�8�Cv�8�U$S6J���N��Q��R��9Ĵ�S�1>c��IO����r�}9g���VE��)�
)w��s:����"�J �h��)������vI�r� �j�u�6	J����U<�����ǠK +�_��aO+�W�Z��=��2�Y)����Ҋa3o�����bY�U~օiSZkqJ�A���Q��,���?̽y��eu-��y����q����8'�q�5vӝ{��5�Y��܌w��$&���N�)��AEE�I��������k�s��{�b��k%��*�����~������'$�^��"�o�J$�L	��=�����410*~p|��zQ&2�q�1�d�	L�L�����L\�᠖���b��o���z�*iK��^뙨Q>c�6\V��8���c�?v\�bT�cO�zLi~ �ׯWNMFj,���W�UT"+ۤ|�����/��rO��꠱��LHijD��x�"�X�* �0ӵ�{�yy|fZ���q� {ҥݙ�p�U��C��|��ޓ�Lib����\�m�I�a�9Q�����7y`�e(-ex��+OL�dJU�ԙ��YIYl��sꌊIv��"/n�t�9�@��;���v}�%����W�81,n�������� O�
V��S49,}H�����x��𪋟��>�|�8{*͇�e����wl������x�>FS�e��M4�d�Zh��E�/\�Id�t05�(\�Bg�d��-V�ߥ���xiY�k=wg�˘oGoA�L��͍^�>���d���8�L(lIm
����i�c�$�Zeo�-C3����}H�s��a^0ϝB�_�n����O��Xʜ�`��kTx���i6�nН|�6�V��v����.��m,w��׭��4�arY�c�ͮ�ǂ$��.li����?�)�W+'ܱ9���b�?@o��+0��(>R�%D�f�A���h6ۨV(��k:��F�*:��+W�Q����4�1R���FZ��=��-ݦ�tWD���b%'�"}�B9�x=ωi�J�V̀J��((��eD���[T3����R 
m���ݟ���#��˾^k�V�u�����}����2{,R����`:XGc������׾�9xՋ�ž��?&(U� �W/F 8�\~�-���\�;�`\Y�|Le��\9��Y��{W1�E3�Zd!W��\�{R�C�C����o�)�!�~���2�jBeZ�]�c�>C;x�N�Ͼ�"<��U,����[��2�Yl�X8�~�Jp�y�Ĺ��a[�C w���_�O_�ߩc4�`8bܤ	�2���Q+�ڌi1�tn��{�@�U���
��V�Jí>6��0u�4s��e���+/ۇ��o��n�*)o�c����[�m�I�&`�8��0���3I�����հ7���G1�Q<Zٿ5��֩�a�c-��"Q5�xSy홭�f��_���dC����x���+o	L��������A�AY<D3�3��դ%`H��X��P�1I����0LH�CTY�mb�v�5��������������>0/�jW��o	9�t�rꩨV�8*6t�^o�GI����>����x2^v���&)��e)y�;�x�Z�I��Yͥ�h-����X���+�Y�6zBU��0��i���T�mK��Q�����:*��+'_�zH\�f�тB Q+���\V�]"��FUa��U�3YO�p��Ș˥K��9�)��� ��'i�D@����'��.�+&�p��hlŌ��?,�>���֌B�n��U�ld�������gVʱ�������[�d�3�9j�GV@�8�C�-!6�K+�R����e�ɵ(S���Fe��B����@��p������=-%�nk�z�,�$���җ8����
�l�����Aa�`��e�������;b�ޣ���4`z�$t�,`��7��S�i�}rT]y�L6�P�m()��ٻ��{hLc���`$L����0`�5���vs$��������C٘���(��rP��[��e��|krL[k
��aO)�5�-D{��ߥ%{%0]h#�CU{���T ���%��u?�XD�3������MYb��e-��CW&��fW�zb'l����3��5.�gͣIQ��[����M	a�Źcg�ܯ��E�t��Uy�5�Q��9Ar����`�>Iļ81���*��P���d�8���\�u�x!^u�s�Z6�D�Ό�t��dT# ��U_:�}⋸⋷bk�¬�E{y��.j4�h�P�F&<GX&�wǙ�����Uk�f3k�S����0�*�-�w�(nF��f��X{�,�E,W��&&,�]6�����5^��J��ޫ��e�l�3��=A�dG�;�@�<Lʅٓ�ކ�FC2j��x���w�b8��]1�Ȱ�~�Ts�	e�4-�P�l�/�w |�|Ū����,�؈+�w�:xO*�s}����O�*�X��1h�wS	F jmAֺ��՘4��f�0�Wkq2Q��W>O��3bP8��{�ef(I���(4��Ia�TV�5Kp9.�]��ʗ�(J�%?+b*In���<�G;%݋s�ؕ���L�i�"o��Wa<.{�m��	���c�VSl�y�6Ԧ���(8�w���F�|��x勞���w&V�fr$0���K��S���qO��}�Z|���qtk�q�������
&55�Z�/����%�����d j9�,����q*�ku0�/!=��LЮ�Q�l�sN�%?�<��=h���V�W캣4����C�h���e�ŅȞ��۔���c ����+q���c[,.a8fL�j���~̵�Mu�cj�2`�q+n��%IƔ=�MT1�b��F��~r�<5V�e�v��9���X�Z���1v�������fOg����o=�W�T�g�N���D��Yh��O)/͏jXٿ��%a2�1#���mί$�"A'��� ��zL�譯�������-�˲�Vp3
Ř;�EɁ�U#K��o3F�X�2i^M�fXVf8��y�y�>����=�49n��$�g�m��e��{2��D�����V�x�>Q��BlS0�R���d��5�7�*�2=�<ݟI�T,��d��
zt�]�_�_��wП6���n��C�������'�;4}֡�� �0Lix��ώ"s�!��!��Е��9���_ڞ��9����9��a����b0��Ky�n`�_�UiG	L����brhT�ca���Tl��t�r�LRYU�9�&����Ll�>�#�&C�������̽)�
i\�;�Ა�w6E��B���vK�*�S#<FL	��wm�'A�D�S�c)�Wz=�sׁ�ϒ?�|ف�0�4����b�������� 4��v��.ίJ�T�1uD�XBd��
+�K]TW�n}n�g�3�d�`�lb���LY<��0��3�p�uR���=�c�����:�4b���=h�g������CޓR/%s�4�c�i�1mx��%2��lG���О��.���d�B�t&�-�j�9���jQ)����F�>������6T�K��`�>&���Y����ؿ6�%佉-U�������?�9���,�4��u<gҷ(6Y2�i�(�����"Zs�nd����
!�'<�[pp�d!��.�4gEc�(�p� �'���{�{]`W⾜�JJw����'h�}��P����II�ԯ;U���^�`:�R/�`�Z�>^���׿g<��t�"gi��M+5�g�������]�#�j��wV��tQ����X��P�^$�F�9��0�"cOp�W;9�R�74)�R���V�a��G;��H��'�N�`+����o�ߥ����SKEp/��:���=�*Kǈ/�h����(�ܓ2ǔ-|N�@�B��ēd�j�	h٦�Q'1>���oR* w��������*��P�Ԕ�( ka^a9\���!�̈-6�R�L��������%@�w�¢�� ����\?:/ܭ3b�3e��̟m
&/^,VV�b����m�:�am�4 H����fV�a���({��MK ZB�T�w��`�#�F<����~�;r�l��V�c4s�Ao�����N𚋟�7��98� ��+������yQɥ�_��8��}��k߾C�`0%�Ag$΁o[-�vP1�Ӽ���g�ˊ���Jt-�G.���=�����Z���L
��� ��5����������*���6��g-�L]�)�сi�O���;��[���TBU5������$�p���K��XM�|�`C�e��4"JLIyŘ��"�H���R���(�9�sL��f���C�t�&��^����$g9�C    IDATX��v�u��[ͷ}b]����������6n�b�~���xB�U�`����槞8z� *�h��ty�>4��e��4��rn�|x��+Y�f$sj�b����^'Ɣ��?���騱�S?zt�
�:�ᅼy�U���T3 �I���<T��6�N8�q��{�ڟz~�ͯĒ��`fKP���1?��Qi+��s)��A7kڶh��`&�4��ȷ��|�����s���o���|��Nrst��&7�~��J����DBXMp�D>�m�`�*j_�Q�S�w����B����6��6sɋ!��9`��h;���FRU+��tB��IW�N���9+��AeFJ2C��l�%�|�f2E�]�5(󑼋FXS����� i��K�Y�$�eJT�ߵT������󖎓	̉ͩ��|�D4�)�#����	FC�Iw���G��н0�쐽�2���,3j������>Rn�)JJ����7��yr\��KW���C)<�&k�+b�93aE��)���R�=��{i�#�(�Dv�!^R�{�`g}Sk}��tO>{�ٷ�aU�g�A�O���[��aξb��R�KƔ=5e#R^>�rP|�f�^�ck�F 0�L6j��0�"���}�:�@��nx����S"I)�	u�ܣ�&I��o� �Ϙ��=�Ñ�)׵��ˮ��n��kFO�+���R|�-��i)�u��B�Ar�_V�~ Pj_������};�~/���B�a��D[fg��&syO��1Q���y)�s#!�5i�k~]������Oez�j�H�u���]�����s��`���/qT"�Jgz�4�'=��TM�ۘ�7��/_�*���c����Kt�6g�\!Y��sVᗎ῿�C����b���PiR��P{JT������T#:�O�%�!�U�Ӌ�y�J��U��8Xޱ�m��;d�\/\�&Hr�9d���&M	��T���,�OqBf F���X,Mc�v�[9f�gmy�*��Э3�d�(ٞc�_X�LPuM��.�}���뇦 ���ő���J|	<ʤ򲸦��������$W�*��hv��Ӓ�8w�bT�w�V�Ņ�#(�(!/��nu���r�8�%Jw�r�e.^p�F��'߃��L
W~T��3����įݢ��S��S&��K@����A�L��x�Q?���k�ם���`��U/�3�;+.e5?��Fq8|�ĕ���>xֆ5���G�T���uS�e�LHY�l��֗� kK��{eL��=�	p���ce�8�"K�b�k��7.Щha����K^�g_�0�3���D�+�bY�X�?�J�/���V~��=�?����Jf��n�/��C��[�Pmİ��Z��3`.� <�'h�H��[YȖ����+h7�bL��u|��)ۦ���U����?(�Sϟı��c)�;k����p{�J�.`�:i�r^�����80��R����֏�h�Q1ƼV��d��$����!ɷ��ɒJ�D�����1%c�'o}�zL)G�y�/I�+90����82m�1�Y���|6�%�
OI����MK|X&�������g6�Sʖl�t����]��׽����ќZA!�zuU��H�x�x�m�,	���="D��^��Y�.��<@�?�J��/���m����>���c�Ǳ��$�����w�`���Y 4��s�S��i?��(:�M1��1��Ȍ!̉Ӿ,��7�$.��q3��$�q
��؁���.����!��C�*��"����\4(�d�:pdt�D��D�}4y�Ñ�Q���%���$_3�&��#��|h$��P�;�0 h��1ˏ�n�rj@���V������0<�'���@��k�{�Qv��x����FR�*�} ��'U`ɀi>j(���� �J ���L"�3�%�v���4�o�O]Wf�=+c3�5q�;�EUkA=�FC�y
(��xU�e��q-Iy��9����kX&cz�S���+�I�B���ڮT�*f�o�ؠ��Z��e4��A����Q��rD���?΁i��������,��l�y����>��O��F��T������͵/z����h�Tt�^5ʙ	�hp�Q��t6���b�H��H�tс~ڋ�c���qeA*��)�M�-]uZ<�Y�lU���G�i�.� %�!��I �/�r�D���ΐ���7Y�ހz�l_�90�4��I#=��n)G�|p��{���\��'�C�	?��ڔ|0��փ��-�EK�(�J'm�Pڸ�HF(��*p���L0��q�����x���ŃN��I"Ϥ�6wM��^�|�������� �t^_Esy?F[5�2�aOץ�����A�[_�6�גn+f�{	?��W�y��3���C�
>�t��	U�T{�!�v�9ޕ����E�%8�(Ε�^9@Y,�EA�[P"Pj.��&D���ؔ���y7O� �� ���Y2��/��YA�y���u}���>-Ck�{���>w�،�ŗ��4��z��AR)�عSE�~��&�+���=䪈�({?p�r{��~��Mbbn�4�e����R����u�T��Y���Ųx�6*&+x��?9���5�y�
�q+�Z�����TO-y������N�ј�����ϻ=��8㔆@)�:ߟ� ��DWT`4n��	\��k��/�{�j]�*-4;{0�,��7��#�3����v�� �y!g�z`��9�[Ͽ}F~��U�4lkR���s�'�8u��|�x���~���ːq��"ُ.��L���K������[Y$�)a�0�{�y���M���#��/|������G9��nǫ�E�l�<���ryw��a��n�b�
ڔ�6�2.b!~�=�4?�K�3�.k\̼Eϛ����%�Tݰǔ�Pk�)zk�9�!�_p�/-�}�f��D�?���\����&��L�1�����ʐ�]݃z�+`���vR�W��h���8b�S&�<��*����$0}��ć�$Y�� �����>�q1������w]�#:�QQ��\�"���\z*�)S^&�|��}�ǔ-l�غ���/�/��ю�PD\�/�cx5��d��Vu��#_��_�gI�������R�2�^q0֦����|�6����>�����P�
��݃Q����h|��O�G�p�@��@9z�֢֫����L�1�p,�%�P����~�!���w�<�҉�֍:����J��7m{���CG��)y��ٽ�HI��v�G0��~�u��|�Ne�� 8�����w5˶@�{uZ4��/\[�u(G>��x	���aB>QV|İ)�L���ݕt��2�`0�0�wh,��X߂��_UȽ����/_b}����J^�/Vn��R�e^�V��9u����
!)���t�vr��Tץm�tH���:�5�W^2�J�US1t.M�W�;!�-�{L�����͏Ę*��L�d~�n��Z4?�ob���5AW�]y����"���lϞ��HFTو�`tb]=���SfFw� �aZa�>d��BŲ�^�{v����:���,=="�ﲂ��4g�	ӹ :�)�w�zNA*��ea#�2��bY��� �k.�u�})3Z�J�
M�7�.}�.�)v8��/���1n@��%+y"��D���(��u�xTU����x�DCuO���爎���4L�w��h����n�g�&�m��p��Dپ-bU��s0�~��0ww�_�q��{)����2�Aq^c���y(^��g቏ܫ����Y�:��*�;�o��w�]���~��>̚��U)�^E�J��ˢ�F��M�W��Iu�h�7���E3�gl���G�"��9� `�0
a�9���5!�3mF�����k5����Pr�R�l`�ڄ��Z���p�߁��S�+٬ZH��9��߇1ius���f�����'K�\��Ƥ�D�[2����"n~�/��]�D��QN���}�����x"�^O/N���p����[vb��E�Jɚ��6ߛ�,.��'��arf�{��e���I��O�.ӣ
�}׌�,L��2�!�(`q�csr��y�eˌ�4v^�A�R^���~X��1
:�Nǘ�0�9�}��}�9x����s2Vh~J�4����2��x�+��M��߹���2&�
2�-�Q�0��fj����<��I�CH�C�v�.��(��U�)w��W���D����٨�����.��,��/�
�W����gGvp�[fJ������L�[��U�i8���#��eW|;-�;�5(�3��S�E�P�qkm���f��:MSZ)2g�	���d�Pl�v]�A�0D��%�Y�n�e*r0���ٷ1�c��:z�7���Qo8��A�1�L���j+q)��i�!�G�jf����c�\+���T$,L�@4��~/�0�ԕ>����\0}���u�?�/1����w�Ώ^���.�.&3d�Q����$�x<q����4�	CC7B�U6@L���1ݹ��_���E6���� b������M�t"S�yjus��A�e�7H,�L}N���\�r��?�}->t��qls.@�w�*V�MO�֐��D�9�˰��_f$@��*���VG��B��wi�/Sͮ�h"gQ9g3�,P;�� ���fW�������D͞��|i��g�մ�1Ie��B���`"��ᄤ�T���P�تFC3����r!������\�d�l.�?Ӏ�bK�QQpU��N5���MTe���l)�wj���+hu;�|u���^O2-6uk��߿�����������K�&����L�g�����v��.y-)3l���ɳGO�}>�-� �.Su�v���p����D�Q�Mgc����рHsL5��-�2p9���b��W޺�C(�ȑ��Y���9ZdL)����-+X�j�w����qu��\2vH���id��N�M]Guj�&{L��Q���x��Q��i�}wҨ��a�
(�07�AFO��g�Rr����\stq�O�0���|�,9��ن�=��W2 у��uy���e\��n�����ZI?&c�a�5����:+ ;�>XV�ӏ&#�@���6%Q.��Lgo
ŗ�T���4c�k0*�x[�i@�~�=�ld�$���s&������/O��-��lO �Ss�u���O�S�`�氧�Z_0����|���}�Ex֏?Z��hb���)U�(�w>v�W񏟾��'bO+�.�ӊ�o��U�"�bU�z~�p�����|	hYm�����X_ ���n��h�Nk?"J�Y\>� �_�g/��o��s�b�u������b�Պ���G5.[.u��I��#����e,��+Zl9A�k%3�>�-1�a�.״2�(SFq�@���8���Mξ� ���}��RJ���*P�����4����{<�m��Ū �9ZAg�|?*���d`��C��.����C���X�F0d�aZ�5�wl׷�W��9u���y~a�#XQϏB�!�:ޱ%�AO#�h�9�YC�6�X�׼�x�S�C�H�?*��z_ �)p����Z|�/��3���?J���TNI�>�v��I ��8#h<��'���5�5[Y$�d�.���JX�1���b��'2Ʀ��k5{j+E�����w��8��'���<�IE������x�wx�������GE��kfq�[�HX�zG�~ ��5Z��5�`2ǈ�x#7�~�1���4P�Q0�6�>�4ǴC`Jg�!�9�t��
��Z��+K�TZjz��+2�6ƴ�n�����}k��+o���,�$���Q���i�67ƴ�Ը�G��ude�pۻ52�j��K��gd���0��Mr^�U����ўn��թ�Ŝw�^S�ڃ�!���U��_���B�q)�ɯB�UJ�B�b�L��g-�Y��0��]1@�[�t��y�0~��ހ׿�Y�v]����l͈bF��5�"�É>K���
cI�P�"���x�N�, ���Fߚ�r��=h���&*X��
�eGLu&ք-D��I�z�Ֆ�5H�AI6e��S�f��qkv�[Q穁��6�D��S�K�ԥ�؈y��Փ���v�;��?0`g��Њf�d�U"��*��f��6�۰����C��C�kn��$�>�'*���#kI{<�,���;�X��_K���x��Kbo�x�w0bD�1�t�2`�5fn��2���Xr�l/ǭXR]"ÒY�G^2����+,�T%*�^�_Cb	��ˣF�i�e"4�8��LR�%Z�����0�~ZIJ\	L۫˚%�>Q�k�vv�l���%�y4��=G5.�E�Ճ�>�$�}~�� [�)`'WJȕ�=�b�F`�-wf�J[:�����
��LW���3�z���
A>�w��מ���8J�]jO�͑0ch��'n������
��j4�cp�P�dn��zF*�^b�-y��Fy�Zbc��-@��H�=��)�Wf��彏N-�FB	t��vX���fa��o��0Xt�*g=�+[�M���ⲃ����b�؋�-e�>�6��/��H�9da���}Eb�d�^մ�9����٘D�"h�om�[xr�0`�z<���h�r|�X�	{�G���ѩ𼧟��=��8�et[�K��s����՛ 7~{S�HW_�=ܷY���*��ɬ"�7�����B������a	2$�v�GR[� f�~}�$i\�e4�"R<��NRa�߱�N���i�:�sߛ��B�E^)׬)��ߝƯXص�<�ǒ� �:��Lj�1����|��ȣ��+��1��X�5��f�3��ƚ�(/Ԗ���B��Jgv
ɵ���a�Wӵd!*����ŭ2ɏ��/b�l���ؕa��iN�6?f�G9+2DS��V�Y�[��.�	�S��]�����*��m�Q����O?�I���p ���pG�f�i����3/x��׾g=��%�P�JEBK�w�|��ѵ-��7݉O}�+��ͷcsXU�iRiK�юd�l����)э�`��gkj�05�H�Z��h\��yy랟YI΀��7�V��y�3*&�c�0@w���~���W.y�k�	�� �N򘾰h�-�2���� >y�͸��_�F��{�nc8�bHI/�$Fe��yRp(G��5U���d졲�]��AUՎ��C���v��M���r�@j}�Zs)�RL��a��	���ָ�����t[c�1ټ�4��nK�&�� �0�R�QGw��:4����u�v��VL�SF�P�t�꤇�x�3���5x�#��h�)�����w����hB����iޞ]�uڱ"��B�s*K���9H�������~���⧪6b�ǝw��w� �;Y�	焙l��:\��`A�[-�,��i��5ya��Lh�A��Ӯ�g>9�V�`��Hx�{���}34�UIy9�Rՠ:�̠�'��l��'�J�L��E�%Ui�1e�eݜ��(k�b��j>&����@W)��`	L}ޜ�<-t���uY����y��c.�ŞZ���97C�e��~���C�\:gb"��6�K-4(k�	TA 8G��Zo��%HoX΀���u�����Zy5d7čI7�K.�~4�hkNi[=ì�伷a�	g�2YqyB�0H�#��([��'`Fa,br��a��q<�И�, Ӕx���E�HJt��4P[���SZV��̽�t$�2K�W�~[+K�lȗ Sc��WX\����఍�a?��Z���3�u�՚ #e)��#��!0u)o�Θ(G��kc��xJ`���dmU���~���WP& ���SJ^,Q���IG=ٱD�SsO��ytPU��[�p�Y���J��F"����TU�,]�eɶ��Ȩ_�N͖�Eb�5�P$�b��*�ΐ��r�*�`�gdd�.X�����Z�v�x�B6T�6���T?�H&3�4%���^����_ ��N��΁~�AF 4\�K0h������Q�1g��~�{+�bD��0!�"��s6A���`>��r���r /������<�,�k���R�AxK㌉̻l��u�    IDAT��'��.��+��2I��S�Z�7,���O���|��>z-q/��_��N�H���Yc�����b�K_�dP\2^YQ,�+��Ql��-_{�~U��BP�����g�����W?==�.�pY�J�;�]��w+[�:��'������e�?��T��*��~3`E�݅+��ّ�ps�l#g�������}�.|z���$L�?��Y��	�dd�9�����u�.Q�D����,(���e�cc]�+�����ɽR�_-HI���7rk�aNE�r�b��hG����V[\x�#��/z:.<�L����Hͨ�ֳ���!M������ʫ����8�>Ƥ���-]wkmi%��%u	~��BN�x�r@�����s
���=�����(�����*ٻֹͯ5�9T��d�F}b�YO��7��x�9�f~���(C��&�7�S����ÿa���{���~_��1[�`g�(��� 3�"2��۔W�NÌc>[��5��9����a����ti�^Ԗ�1%0Uδ�Ǵ
Ɂ��K
�y�8�;
���h6�'���\�9�U`�c#kL�0���(�=dL���TĘFK��qI�}J �6!�'.�:��1���������Iy�ٜ���n�;>|�zLG�%��T�5�
�g�(��u���i�d��J��5*���BLg�5��G�����xً�7)�'[�����e��Y>rB̕��~�Kj����4���U3&���K����A+g�QU�M4��!l�ϚMР�{>�������\���2��p�Ȁ=���}���M4�a��}hrl��������|�	���4+��{ܚ1�9��*�L�n�h�!e��S�[�<1 ����J�)�-��v*�LlJȰ\x�?C��H�������kQ���ԥ��!��\39�R:�F�Ik{�{�2�F�QQ���e֚�`�3 �"���s�D�[ OɅ;�M�k�&,�i�#��9tV:h4�`gI=�� 7@ȿ�����6S"6��$_6`�	���2ّ�c�S�=đ��_DE=�����YV�ӑ�*�ဨ���'ב��~qF�W��!����,��Yܫ�T9~uI���بwWA� {��, �L��������t&�:
J�5.f7cZA�}[L'[;L9�l���L�k�iȾ̨�lhE��R�bm��XIRg�m���%�&(��h�ܕs6�S�IeoU S?l2]��}���!�ܷhVO{s�vI�g�)f�$<e�s������O�キ�%��3�1�=�M�Yw%riM�z�����90��,��׽�}/~��LO�m���x�
d�?LrM����]x+�����ꃶ�K���_��T��?���鮤(����u��u��l��4���n �ݣ�ԾZ2I��R�1De��|����^���?�,<�&:n�kZf{>�� us|�m\������
6�uT���^ޯ��y�L��m�sy�q�[�ï��[�ѸG���bO4+R,<��i$6~�3�N�;U��`^	�0��l�K6���+9������n�*�����d�v��+�K[!u�%��1<�=��3/֩�v6�3z�X�>�
�*��V�u5����-�4P�ޭІ�n��u�!W�.{��1�����5f�>b^�124�'i�2����~��ӹ�{;ZE�ņ��|ښ�i���l����y�aWgV^����l�2���-��}T�u��������t�-S:X-���u�g+�����_����:����csPŴ��^(T]L�t�m��j�^��/
e�6�!WQ�O`�?�����޵c۴�L"�$R2'��-)���D2��z�i��mM�T���g=oz�ph���3/�]!����[s�к�O?y�qٕ7��9�cPXc��L�_�4�mkݶ�ܴ�S[C|�-�iIq���g%0���6VW1k�8�LT�kSc�ve�PQ����ɘJ��mb<�h�]����h�е��J��q��9�R1��1�K�#s啢��vY�Q,�|k��=�4�$0�x���\���z<����u`�����.���qx���ҡ��{���f��LghT��$� '�}.\���`=\�9�3i�0�>��p݇?��_�K���8p��OlN��^\��p�غ L�J@:c*�uV;+s�z�!<�IO�c�y��7��-\���`mm��Ih�z-�tku����TS����lb�����W����t	^���ɀ��q\��� x����{��9^�o������ù#HK)'b��ˠ�W�����LӑV��*y���&�c�Y�$ؘ��2��cRǥDa E����E@��V&_���N���XJ7B�h��>F#UтM�I,�p:T�5�	��:�@렣!�t���F��dn��L�a�Y����Uճ#�G���$ћգ�����k�?��L6�v>g:�5���]�J�MH�#S��b�B��CR=�9�roJ��+�
��B^A�!f��6�h�;��ʓwKq��5������98ex�z��XkNm0��F��|bCc'?��N@	d#��;C��W�0o�l-��pPj̊����p���߃����a�CX9xH����0q����&@�(08��9�z��
�4h;0V8��nA���TS^+��뛨��tH	m݆�k��z]�R�d��d���l���2�2��Ί\�<\j,h�& �DFc�Y.�H	_���+��eLg��(Ō�,���;����`s7�X�����@�}��T���(�EcG���tӾ�ّlMck�:�����ؤ^���&��Lⓣ��;�ʞ�{�D&��U2�C2g��B����%a2��)��pپqӣ�yz0L��NE����@�$|������
���w�S�7P��G�X�9?�7�̋p��g��Ѻ����-��8C�[ �޸��|�r���#�U1�u0�4�j�V���۫ gE8L4��NT1��V,�3�4 
�i��`�����L�L�&8%�,��db��b����p��3�m����ޑ��}�k2�����W^ P��,\g\H��@�Ai�eV�������%M�+�CF�j��x��0�����s�#n�{è0}�F�˳}��=�؞�k�O)�\���ᅁ|_:d�
���(�#RJ�--�������v�{�k`��$KtOk;��Q��8�ӳ,�'��s���p�8��s�!<�O���;}���!q1�������p�m\����图��7�����.
2q�&:˫�ͫO,ۊ��0+,��|�A�U�%
ݱ�e��4ªR� UQ�ol^�n�-F�r2�^���^��ç=4�<�3K�����4�S���t��R�{������)�#��R���f�����{?�Y�vw�bg�9���aƎ�f˦o0�贁��-�K�I`Z7�t������z<G�)Z�+h���N���O�:� �:Պ1��\y��c�G�j^ L[��@�E�����w�%�U�)U^��=��kd��Q8�2�����y��D�XL�-���1��?0���g�czO8.f�4�jⵀ;?�ao�Iu��ӘQU���,H�f�c�[��)�o�l@`z�����z޹�1�����g��ݸ��/b�3В8�o	++m�]]A�f5�6N>t �|���'=��rP��n��p͗p�wck��q1�`4�����;E�N�`:�KjAƴ�>�k�Ϳ�F���g�E�\�cT�
��������x#����٪c��)S�R�al�_�U���tY�=�"*�ـ�z�N-VR�!Q���6h͉O��B�&^�ҁL�$x,A��>��1Ӧ��)_�ou	vF�A������2���L�϶���vI�(s�L���r�n����L)�6Yd0�C�o.f�3��U�w��B|<�J��I<ן*9.�B& >��Z~p��f��f����j�e���+���:N��Y�J㐣Y���J��΀�sc8��u���%�/Kf�7��ˣ��?2wP�ΦJ�`F
�Y?���3�찥�!��J�[��K�9�l" X��cJv�8�Bå�g���Z������U�i �e�n$�b�I�m&$�I5s��d}ӭ�~�y6V��ڿ_3T	L94�Uf�"z�{�j���@f0�d}K�-S1 2G�wF��L����6�,PZhFi�#�����*�9c�	�1P
�pzTi�%Gr�رW5U�����n��#�����f�&�LR�_[<{��2W^K�?�fic��*�g�^bQw%y2�6����Y���ܔ}1�����Z�� ��e�8�ڌVStX��,Q��%��)fw������h��{������߸��g�����43����z�'�X�i�w��'6:�As�u���zO5��33�(��c>\ǩ{�x�3���^�T�}�^,c�;7�����j?�{��q��wpٕ��[c{�D��S4�Pq�t�Ӕ7 G�	@����'w$5���lU5��$E��>;�<�:G)7s۲0a�B����t�\6�x��i���Xo�?I��\;F���2�k����j�rO�z��̙L�����k-XĴG���=?�cr60R�T�R��aV���%|���v��G�J.KL�k�V�"�B@j!Q��+(bq��i�b�WQ�-{B݌S���,���F���^鰜 V*gq>ŤX����m�G6v�m*y�T�!�;'М�ph��g��H�'>f��v�lYl�'�m��O�����3�ބ+�����qL�+(�D�sI�GZ�6T��1�ɦ���Aۋ���X��oJ������sXS�I�����gH��F\�ň��Q�jD��S�����ڵ.x�x�/�g��vSKS��,������gkk0k��J=!u\?8:�/�
��t7�:��F��"$��B7Z�_���fS��LY@��v��Qv��-7�1/�T�`P�B )oˁ)��TԄ��l*W�.j�i�N`z�����r�_� ��4��M��mj�)��u���(�1��	�f+�(/�j�.ϋ��
����i��Ms��O��h�b�v��÷�O}��o������jL���h~-�Hr$M�e��V3@"Cj�GƞVg��P�D�#��ş��/�'/z�B��=����w~ W]}=:�&.|ʏ�i<	OZ��ʒ���v��n��f��F�d�?(0�0&���O��������o�UW߀��]W/[�]�d������_z^�ܧ�ݰx�9�}��}��7���:�/֍��rA�����̯�Y��@1A���R�pv�c(�S4:�;�Ro2��T��b@v��vb�%N�G��8ɔ���%8v�9R����}��'���HӢJ��FQǮ�5�!)5�d�9\fA�rd�87�f�&�h��%}�2@WѤ�j��Ʉ2m&��a��`& �IIA�Ϥ�$��*�(YQ�o��y2;
�^E��A��S�7&�^1g��'{�CF���1�l��Vd�(ta�i8�R*��K@ቋ��BB�d;ˣ���>??���v���d^��|]�A^�0�nɜ�S���q�3�^s��ݐP��G*<(�6�"9����zL��फS%�|L�'�t����;t2�,k�$�>bo[U�)��)�^��lۀ)�z}y	݃'�����:�X��RP�@`Ze�� ��0�ؖ����7I�-K�� �4e�bK�(��ɽ�,�4�a�d�� x�W��~�a�a΢����X.%��|L&gX��R�E� c��e�%�fG2��1�es�b��%CI�d?ߌR���,�5���h)7�g�	�m�ދw錙g�)q�G�H���k#11���d�\�e�%X��bX��$;�ȶ��޳\'=�u�Ec���+�=�ր��+���U�����E(��lIa����u���Hq��1�[[��}[�!&�-��h���>� ^���yO2N�_�!���.:�D�#��'5�w�;�e��>q�������˨4hT�2eO�ZN؊1��^X���)^>-��J��/ӄr]�f`ѯdA,x��,
��i@{��;�Gq`�������CUl�������;TGO�K�n�w����@9�e �(2Ǿ�-�1hS�CV��T.�t-b_3�2�WrC.�]r��{���e�v����D &]W����Qc�amD�/bF܃@�� ��`�j�}V�Hr�h�I3c����
gvq/q]q�����\�"� �~�Q��oWFX�q��������Sp�~����Y&���^E�1���n�����ڷ��	���2����Tv�Ф�=c�r����z���L�Z�QT�3`oaԞI�����Hs�-�Yh�,�e�ސ:�ߔ+y��F`�͘`��R�Щn���_�"�g��ǦT�XX��(ϚhGH�Eih[�ӟ�	ҍ��]���3�6l�3�F�.�4�lT�_��y�7��|�90���hk!���{����֢�
��첽�0�t�#Z���[��6�i��R���ӄ�2��Y|�ɕwO�=�L�cz�a}���&V�N�LELp�Y(8��Ulf��笜C��0Du�Ge��S����7�,���SL����_ɕ�#��� cZ�1j���ҕ�zxBצb3�	���L",'�3`*A��d����騇��1�jq�/z��+/��o���A��[�ȳ��Ͻ�x�cd��ǳ�-ĞJ��8�H)@�|�O�V|�×�{߾����Ý�8�P��k����/��<�3�����8r�@�U�I�NB�CsP������f���&�rPJ	�zv�_��o�dþ2���E���hδ�����p��s�X�f�	��J��Q����x�S�Q�3p&���픽�LPFF����J:���ڂcRƀ��?gY� �F!U�ɕ��ʑuc&�gK@P��bG�!�X"muc����Y��j6Z�G6O�=�C��
��d"��qV�{����n.ut��4"��qM~l��D���A���Z�ze�-�t�c�fFԜ����̘ˁ���Q�0Y�'�b|��*}�˅�IE��$�fB�+K�\��z��DN]�ڷ��;(�-I���#fah�+pJ	�zDe(UZ��T��Z��y�Ŭ�9�;�d,���j�T�,н��G\��d)����xsK,;G�4VV�=x ӑfk�hk�+A[K�\o�d�d;���X��+HE�H����a-1�-�4Sv����ݚɎ�}xJ���
��a[qʐ�ɫ<a���k��A��V�"��X$}!/s��U��5�z��胸=CG�H��gX���9�:Xl���Pv�d �z��}K0��/�OF_�V) �>��ђ�	0��ț_j�(�9ѥ�/����ڸ������R�ck���gJ��!.�"�p��љhŦ��7R���W*�y����ޟ��[?��b��JŹ�M2�g��1�9���Q,7&8�qg�׽Ox��Xf��^35
V$���Wm�����{��ا��O}�Fݜ��ڏj��z�+�3���&��ҩ�I��#
hz�vgR	Xm��Q�=��!�O��� מo�L��ҞpDz�.u�4A^zs
��Ou멅�L&����s�u�O�*�eδL�u6{�����@P����{�Vn�k�i�,��y?ik�I��ڨb:B����qi�%��?,�T��,pg�BY�yP��5��5Y�.���>�����m5��s�/��E�k_��IrŋzI!�:�w�B��L�Ln.������-TkLFr�~��p�k^��x�~�M��T؈�l�;�YNzl��go�/��}M,i���z�͗�Y�fL�v��0,����(�e�(�����t�2�	��
��C��y��\�%󎉽j-+ڲ�A�����w}4�C{~���^��{�S�uAE�����������(�/����R�{��M���7}�>l��Nk(fs�n�Ui���ΚL�K�7���z]��^_��lD ���D
.2��~m��S_�̕i���l�F��l_C��+�E�t�^Ժ�$���Q �&�uL�?r��P�$�p���C��U������7Lɘr4���jMШv60�`����k�'��6��0wN(    IDAT��+��|NWޏ^}�ꃟ����y��Ua�L��%H@��'/�8����L#bX-���3 iD�q_�t>�D}z�����>�1R޻���_����f���G�?���p��K6p8�:�B-�P�	��"�ܡt�D����\����}LF��t�������z�𬧟��[��r�黮�>v��O�1=t��|$�M�d5�1/���61�D��EI�b>g�ɪrF"�i�����:w�t��/��9	v���j���,PJ��@��F���t�<�V��UQ�72��
s8��b<D1�Sr�]͘�#,�f�m�L0|��J7em��L�����R:$�0%��h
D���q��M�jsA�[H��$ǌ�Fz���a�9#�eCv�P���tn ����X��4k�˶b�1��{��T�<�j4�m)��J�n����������*�U�e���^	2RҞ�˔����u�	R8�P��H$OO����g^-��mq���dЌyw�Uև���]�/R���X���ʀh��i�f~���wVY6`J)�ۇ�+/�U��cZq`��g��P�&i��ol��ّ�����*�����Ƹ��	���8(�2�O�{�o�Pc5��^H�K3��p�%�{A��2�I���'�d�U�\u^�"�#a�+��f�6�D��)�pbr2� <A�g{�ΙMϭ�2J$�H�5'��g�މ>����.��~'=�I��������y���]�u!3wW�(�(-YG�TD��`�u����f��:����sp.�5�F;�Nn���ᅟ��כ�]@!�_�X���QXv�VPJ�x�sb?�����ZT ����bT��E����Ȣ�f+�i�|��p�ͣmþ�?y�S��?�9�TT;C���L>�̃ u�|��M��#W��܃^Qǘ^��6�<�8$���%�����+�x<U!������P��3���Y�ƚ���3�4ںq�Y�EL����s��b�}�ֿ�S�0��?��iXH\��y�ƶ9x�����fs�p_��,fm�"j�}�����auUF ��@j�Tʓ���q��z���A�� ,!U�/��;�.�G���7����o���/��1N]{��U����be�7���\_��P̚WdSxm��㴓�p�s_t�>b�ؚ�&���}����F��7� ���p�׾��QE��J}	��j4�l4�];�#�)�vS{�)﵄��P=׮�pU�Σ𧈂_>�ܺ�J~;�m�G8�Gnn]�,*M�r�2^̆ha���ޯ�oxΓ��R�o����'���gh�L���?���<���vl���Mw.7tJaѢ/�&u�G7#Eu+T+hҋ�^S�Ҽ7P��ll*@cLWQ�.aN�I)��*S����)s�L$��/-���̗��'�t�0W�ɕ��G�1���+��nkj���^؈g�����	L�3aΎ7Ɣ������x��O�&�3�L/�����~GgL'��%���6�U���r������S2�59dV�!�2?�0�o�f<�i��щ�H�{7�o7�y�wp�y��%o�<�!��b��}qج�r�u��&vl�����\��_�]5�v����Q?	���7�����'+cTL����
���8�9���С�:��[:�b���Ƭ��{�h�F�q�����K�9Vdշ˄�,"+�d�<ٝ_^�jl˚��X��`�1�5��=E���ZkI U}�~���/{)���Q�a8����9+}�hVGؿ��2��X$+E�ө��}�a@�8;��k	)�Yll��Z�K2���3��8�9��9�x_�mڬ+Q�hfR@w�|���Oq9�E��uTf#�_��p����d)����T:����J�dJ��ϰw�M�Y�d@+tPk��z ���u9��ߝP�
�=|�K����CS	[0�:Aʑr��*o8Wz�`��p�;���gɬ��� qwLVys�l��j�m�F�<=������It�n�,(� H�S>cЯ� Ӏ�ۇ��1eP�{蠀�`��Ô�`��ߌ����tBF�����=+
����ɎW]^�g�q3u��>f;bL)V"#nx��s��R[3Ky��4��k2tK���8��oV9C�CIwYX��#Y����L=w�7���(-Nk�N�ZTf{�A���J�w��%��3"�޻�dK���=X�c
�t�F��b^��Ѕ�(d��&E2m�LOJ�m??*�Z�N��=�!��OK��i�׾�����z�ʔ>��<�̿ln���$�,��}�ޓKu�q����6ƣ����_������{��y��m�Nٻ�IXƟԸq�#�O`��=2|�#O�O��x�3��i�:raT*���'�޷\���㊫o�U_��Y�{mI�4�k���9~-�]�\�h�4�*ǂɍ���;��J_q���Br,�;��#��������x��?�?� �{.�*>gS�iw�Fӥ�����J�|���L�
2����y�݅�I;���ʟ�Zw��J�����X����7V�u$����[|�90M�a�z�k�V��54��ŢZ*�\�d��|
�Q�<�> ��O�bW�o��9N.m��07�cYS�E� 0�l<���ơ=5<�)g���_���9'��a_�����l4vL��3������7���j�r�qLj+�����誏4Fۑ)�F�s���zn�)ђS��.�*,����?Q�z���(�Xˊ�א���J_�MH��SW#����F�s�x��Z�-�}r�;��35��U������y�&bO�tU�p�����������;l+Lh	�o+�/%k��`ڨi�A0��8�À�\�J�3�I��L&&��vAWV�5o��e�Z�X�����y;k�_������{��Ϧ'H S�����<i:�đ�0�јt&㦕}�P�3-��X��T�2����	���M���2�:�ĩ�~�W_#`�����!0��ڻL�/�_�bC�;`�"<�dc�>aBcjA�� 8����&�)���	�ƛ�M�����-x�S�
� w޳�������7��X\�W�ag���R��ɰ�,,_�־����m��k���?|%���r�]��Шp�ه��o��w�W�m�瘒1������f���5�J3.Ǩ����g>	?�ܧ`�2�TL�ө%;ƒ�f����Uec���i/�@���Ȟ�Q�*�o}����]|���1(�Ƞ
�9sX�WafL�l�'?�x���!��þ�%�SE�3�i�7Peˮ98c,��5��w����3���w���x��v_��V�u�浖�$�2���\1�@l�x�g�&��+-���Gࡧ�j��ev6J�޹�k�+�2 #�MN�x�*�1��N$�Qy���1�ΰ�=�]�7�N`g\Ŕ�T���P?%�mVdvYQ�.���JP�&W��+�y�Z<�<a�=�7�:��Ε�4�<=�)Iɳ c(�J��GY�+���ݮXS�*\��DRnؠ;z]s<	L��L+�w�!��|#��<`��"�]��!��m`�H�;�L.u�{L��5x�,�C&1���O�ţ�>��c�ے��RFwܝ��2RJ�H0]L�L�Ԡ��[jX����
*b�lS0�!���2��T��H�cD?K���c�&㕒)�D˝�C�	�Y���'ә� }���D��-���j��`?����S��u�NFi.���ٺ�������*�����#��G���?�#92�����P����V�����T�*��,�n6�ؾ.�VO�+,�3�>�'A����Y���:##�0��F�Ě����go:�Do�^t�\p��ꟾOy�#������G){/%Ӄ)p�1��߆�>����;��=F1����N���
ڝ%4-��>��t��A�#�\/�\���z��(�NLYЯ�B���@0�Ώ	�]�����Z?¿�4�B��
�����J�`�����)o��D�������U�#,x�1aMk�G܏�I�q��~����6bE^L�u�ǲ�am�D��癮�94�ǅ�]	ҍ
\��w����@'PgquN��CTY��B	��ڦ����NF���b�*n�C��xʓ�g=��8�1���Sk2��n�q����\����z�]y���Vܷ5�Lka�,C#�FDa�JMf�ǳ*��T�E����ޕ_��i�J��(`��������S���k����2�z���A����Ae�Cw���?�,���ހ����q�����vĿǿ��l.�`��	|�W�򫾁�6�U��SlH#cJ7^���0���L� i�%c=���M2y6�St��0���a��ĵJb��K�]��+�;�N`:�_J̀�>3?ba�^e�&c�G�cʶ�G�I����vK�G�e��nvB6�Qj&�%0�bVP�X �dL��O��X�׀i�R�K������I���$��T�5��tҥ�a�`��XȽl��H�EU�"�6��1m������6<낳cJ`z���ӷ�=n�廸����_�2����c	9�-,��V��1��r��ͱp��n�>|%�z�70N��TG�:��9���KpޓNO���TR޿�<>�����M]�سg��Fm��l��Z��+?��>�Tt�����yX ���p_�Lb�J�
��Hz�<bQ���C�@��4�W}�������Ļ�����L*��M0f�mb�R�?����cZ��pY��ǤE�)�3S�����C�-XR���1�r�pl�����{>��m�1(�[h�h0m6Qb\Pb����I������g��TտLn�����]��o�
��t/�/�9KH�� ҟ ������1|��GQT����;�@U�+J��pb@Y�E��)��(���'
.�kc~�-ʽ�е��vX�P��:��p���>]�����V���3�H�;����\.v1����Aޤ���t�i�b�J������ؙd)t����a2�Q5��h��蚔��~�b	4�\Vr*����c��#S"�F�D�L��){�:�v[��������svC63�E����1��t����1�WJ�|��ܨ,6W΢g .��A�B�
�Yb&��_��X�+��A=q2-��R�l��cY��J��	��{p
�+���zC�s�Z���Rumc�r	�Cƒ
�m�)���|����:�9��S�U��2�R�̓9	��V&n|���E�EF®��x��'��Z����<[�H���3� �gH�B�HIu�Ş�t��"�x�c�xa1B�>��b�]���y
^����a��A�(6�f�'�1Ι)pt����w����F��c�XB{e?�K��tV��p4��l�1�*xhOQ�W�CBj����`��<7�F��;+]Z����o��=��s|eF .+��ț(���^4
��Iѭ7��.I�[.�X�L��Q�7`��S�#��$�q�Z�a<������ S�;e�RLP �X�`0-=7���pf�������(^SZc��i������	|�r��E`�Jf�Q~��؈���t����J2`BB���(t�p��lBs�M��}X���?�x�ExܣN��ղ�������cD͍�y�1|��W�K7ݎ�>0o�q�sHk��;R�՛-�#�i����7l�]�+
$�7�ܦ�v�m�W�Q!��P����=,v9/[q���aJ/�8SjY���,�$�`�������/�k~�|����a_��!��
1٭��gY�*	�Xa�k�� ���+���^�E;�)8W�#^ȖV��1�\tK3у1m�E��k����u)�h�:����}��fS�|1�����c:׸�.[-(_���-54�Kh�]5�#���K�լs��4��l��q��Q�1�zJy��c>����!��b�T�'^��Ѵ/�4�ǝ")/s��1)���|>�1��N��{?�#��e���:왩s������+�yP�qe�)es����T՘[)��߇I�:�m�ş����G,0�wܽ�����·�u���^�<���A�IuS��򬅀K�U/��k5�މ���Ӹ�o`6�b��@m��{�zL	L��Uu�����|貛p|s�N�c�tZ�Y���k�;o}�z�6�|�v�����L-�$ �h�v {{�'eV�qF�g������'�k�6���]B��mo?I�C��&��@��<�!�����8mժ-Òz���߅�2軓[�D���\�I?]QU;P��ފA��������4�y�	��54�-t���Ƅ�ЩV�p��͍㘍���=�+~��x��^���ZP˄�V	6bW�B<�x���sF��EAA놃�࿿�*\z�W1�������)�7��a�ao}�Q��w��-;���-����^�D�������N.��/u�ngY��ޫ�]�C�$�� ��ۨc�qfP��RGř��`����b�"�"-CMB��{�^�u?������9�9�?s2I��^�[�������}?�#�����BÂ��¯Oq��[u�D�it�%f~D�ڤ�����\E棽t¨	c�B��@� ��㲰ɘ.��;뵠I?�Hp�Z�`\Lel�*��6h���Gj�_�Fh��g�|l)O����c��1-��b���k�%Jy�ү�(��C&�1B�>�N��6iTPE}�, Zz��ȤzM�����:���פ�'	s�\�35Ӳ��oQ�Ʉ��\���:��=�0���̕�ςBX��}���2�6�8gL}����F5���2�<ѽ������qD���2uֻ�`����H�l��釞�5�m�Ē>7{�b�U���`�_ALP ��@fi�Gf�$��|xc�]�i���luf�8;�z�{�`���fq�!�2�taQX�N��iBB���*��*�`�Q���z!N]�
��e%Q��Ѷ.��bb�c�&@��7o�n��w=���&�,"[F,�C:STQ2~f�p�ğg'��'�I�ٲw�3r&��k��iϡ`�AU�1)��VY������iQ¥璄��<����� l����f3>�6�WH{����Lö�v#v����&�u���3��u~~?�-�L��{��@�]����^���	u��}�� �e���f-����7���#�� mP�,��3+��ߋ�$���Ф�b��%�ji�'pҺ�q�	+��O�� #6�:dHuo۪U��"�#ݹ{wݿ���xd�$fZYtS�@J�h.߇nW�dY���hs}͝�?��Z�	Z��9��^�%�9��TU�l��5gT��Q�8�ϖN�^ؐ�3Aց׈���p[F��+��m8k�����$���`�� `����6a��`:]'c�`�e��e���q�����$���b��c2}��^��Vg�ѯ=��LZ��R8�KXS3��KgDeV���ظ0�,���y$��?��3�WUO%�L�9�$�`:~�ꥪ��LC�cJe�����B'f�3�*�dF��W�v��G`:��}m|�]��3�-��͏B��q|�{7��J<��4$�6���>�v���h�ey3�TI�6Æ,��_L�ݸ �n�.��]E!Q��/�g?�����c���N۰oz�˱v�:����è�"��m�u�VC�^C�V�}�l7ݵ�����㦻�f3�&X��\t�98e�b:4z��|�k���f+�g螜��`�l�t��x���s����o��k登0;G���ŭ���:"��aM��1��{2�1���	\��_¡��A���H���Rν�K�i����lBO�&�K��Ct����b^}�8$��+t���>-�F<9��i��2T��{�|��q���hu9� �\>'���˲H2�j���уh�qz ����%x�kOG����wK^t�o��	N��8LE$g��ES�_;`x�3��o�W�{#��a�b��ugļJe�&9�qa����P�#�B������*��r�hba�P[K�uΠ�0���������b    IDAT*�9���D;bã"\�bp��?�K��8���'��z�P��+�4�hi��؄ē�ysѿx!�26I}c���~�)�A�შ�P��B�R�bX�ٰ��C��j~d=��X�+����F[y[�%ěz(�����.ڜ�HPJ<E��V�g�i��.2����И.IO�dAE�	�9��D$��uɵ#��r;a��M��� 9����m�����me���Y�SB�*���ѓ�@F�.�
y7qұ�y��aQ$��Ä�gK�{��.(���q��0�M��� m�{�l�8X̮ޯ �c��N�����
@��{�34�������ls�:�%ﳍ��g�0��'�����x�X`\$֒��rssF*�:{��hW'kLa0�=v9��ux�'bn��S�Q�T��k*_��C�?�8��aܼq�3�F'�dz�l?2��2nF�i�f�ztcLo�����Wf�"ʓ@5�Q5���<{q9�y`�d�}��Zj��˂�|�y� 7��/�U	>#&m��	AU4f*�����b���I�DP�=�V��KL^�>�?�#?-���`��Q.�@a�ņsCU�kϝ�%������
s<����OE�Z1-��e}�AP��.ٗT$�F�Ϩ~=.M֢��-�:�	���������� R��4��2�*2�&�;j�>}^��3q̊,�:1I[N�]� c�H���M���{�[�G���%[�E;�G7��.}6X�##�<m[�����H�Ӹ2�a>-(�P�>�0Kү��=Gv�==t!��,�:G�+����N�S�E��V��X��*H�𥏿동#�G:l�ڍ��3��'�˗�0�k�{���on�?��F��S���0Y�L;�n2���\�\MS�e�}K��c%��\��2��Ҷ�׮w�H��!V�ƕ?�7�?=jD�ۍ��Y��C�(OL�Y#��mW���ɡ.��:��k��s.�b&��L	����Z,�S�.��:'�S��bĥ�~��F��că� =@¿:b�2������ݯ���f~txD�h{80�ӼX�3yf�I��6�z���0 ��0�lʵ�JA���7�8��j5�(孎	0����S�����U_�6޹[����e8���(57�{X-&�L���)LMM	P��;�n�ķ��5n�ݝ�ֺLӉ֯[���G�|�B�|�l�+������1^�BJ`��˦�6��
��M���V́�вK����&����4�5�9̟7Wi�Y�ɏ}�z��,B>E3������[�q��q �����0�$r����r�T��iHb�jO�eg��e�����G�P�Y_������z?}!�!�?~D��!�>���q_��t����̵�ş��n�|?��l L��өʥ)L���VŢ�$��߽oz�i��z�@�tD�%KDTBn)Ch������2ĒǙ�
ͣ�����p���G#6,s�R�"��5���>q	
[,� �GzX�k�|k&e�9֮�=��ϊ�=����碲$�z��wW��GF�7��{�&ɲ���A�lf,{I�
��mM��p�Lq���g��@�zLy�b~�p>	z���?A>;�~2^tcRA�U��4��>c7B����A��ƶe��!# w�zK�i{���G�M4�zL���#�4ƙ���Ƙ���0Ip����?�l�JU������C\V�%~*U�b;ef���?�MF_j�-L���I���_�+�o�Ji g���[b��,�4��d�yq�.Gס&B���dLS	aK ��X��,�غ7��VŅZ�,[��}��蝞m��Č��݂���>O����A�sh��
r�q�Ẕ�7���H���%���tK���lHȀ���m�\�y��dm�s+]z,�W�F\9�{�4�F	�n��8r�6�^�W��9b��O��5�����H��]t�
��[�mw>���عk��NH��Rp��HH-ʸ�X�=s:�������Q�Ocƀ�\^&l朮���u!��uM�e0�!��~r����0���&;� �%��:�'��$�k��տ�bF
[�&}��@��S�z����������g�D��=h7����{�?=��Z�!+0�3��}A�[���R�m%R�+�^���m�]�T =��}�L�X��xm���̇�6��4�aѪ��m�ѩM�?lX�/z�8����lQst?����j-��ӄ����w㏷ߍ��/�]�;1�襐�d?P�N_-���j��"'���We��%"��^l�][��
%�ح������z��g��P?]�X��g^���A���?�
9�4֩ +aN��k���-�3��0��9������;��g�Ԩ����
0=4��t�6�l�L�/�-�Сy�S�f��TSR2�i2�3%Ԍ1��c?h���X_?Z��3"�+I���%���qT&gЬӸ��L���@?R}��ʜ��N����Q9�C��8�*�	L+U�w`:�n*����Z�G�=v^��(�8�6'�0W�'.x3�8~�Hy���kx��m�	cJ)o5Ι5�����֯&��kD*$����F��S����9�[�J�i�:��T_���x�I+`�ͽ��|���bǎGq�'⍯y)�]9_z:��İ����j47�T�R�9��'�e�t��1|�?�Ϳ݄X#&��L��O\����8y�B�_4'��U_���݃��"�M��Wil*іJ��!�_/�[qf���.Y�v���x��P�T�����#W��O�@�%D~�8���Չ�����{�!��ahhs���KQ�i��G��b�y�'��H��|��5�d�G��Y�7�7��W�^�y�k�Os`�}Z�D�	�ٻ{��G�\F__G�X�yÃ23OM��EW �	*�htQ����@&�D&Ê��8&��m�N�k~�M��A���%&-��gş�u�^�`rb��X�ǹ�J��է��m�~ w�bv293���Q̔�X��x䳄5a������2v�ُn<�X<%�K2�&C.��^�\.��NB�����>v�q2�E�r}b��M�dD����6�r�'�>�ð�*��[΂ȚA�H��"L>f�Xg�����s9��u�AS���i>�M�CK�t$LW䮉]�2�z
�h*~f�:�-��F�������o��C+I�^`*@�rD�qd]y'���V�MM`g�O%Ay���PVZ� o��j�1��oq����5m"cJ`�/��J
X��bA��]a��_V09�nd��E6�9b��^?^lP�g5��?I�,�d�5����GA�0��0.I���@Nf`%ܺ�$�9�����*G��G����L�d����j5)/�$:�l�Z�����n�aV�B-ɒ��OEϧ{Ӆ��g��m����"���<e�d���cN���dg�-��������'������^� �|f�M�(�=�Qa����i�l�?�`��J�����%��4y�D��_�׿�E8m�J�%�jn��=W���ߏ?	��W����܌Gw��T�D�d�t��d����i$�4�S�%`�����Q^�.���.�-�ɹ����q`ʘ,�� QtM̫7em���{����x�������R�P��a�N��g�*+=tok�@W���:�C�O�����a=�q�^���N{g��O����r���)�)蔳�
��G�U�'{�#_ӃG���Y�C�xg���8����F����&�aUOh���i8��֭Z��j�	dbu�b>�8�x�u���p�Y�����9$�6�\̼ �Ľ�;Tǟ�}?���xl��bĐG��?��op�����PŃ��ʩ�FT��~���]%`�r�"$�wnl\�_��j���@�,`��]SR��)��w��>%ɑ��:b�2��i�����+ߏUK
�P��?�F�Á���'�����w�ď~~�Ot12��x�F�txR`�B-�K"�5�f+���a��f�̀��e>n�i�Pԟ�n�^&����8��$ҭJ��LϠUgG)���"�Y����Ԛ-��AU+.y�TZ�F���5+̤��)��dAQ���MQ���.��7{Lu�)���TW^zN[5WF*9��d����=�?� �Z��w��.Z���X�#ƚ�iV�?���M ���f|čC���7�^Cmr���/Y�W>�A��nIp�<�v=A��;xh�#x�)���W�Ǔ1M*�'UM�%j�>�(��~Z�8�
Rʻi�������4b��N���dLOXHy9�����k~�_��!�����س٩!�-c���������-P���b�T�u��>/=�s��%��G_��L:eFA���:c���v��+��ǟ����ǭ�{�q���2Hz��ۦ��f�08w�<7����V��UtZ��x�������l�Ul����;��|�\��	k��IND1������P$���S]n߸7��6��O"�J��u��5�y�Ō$�|dy��ħ��%6߿�V�� �}t�S`�	�)T1r� J�x(�����𺗝�>V�-�1qܺu�?� v��)��o}�[�W��㉳
0y|~}�M�?6���
���/��:���<�-]�<�Y8��c�a5���{Fq��?�F|.Z�"��2t�Q7\q��5�H"�IO_i40�~�Y�H�	��Y8L��o�x�F%���a�B���7�}ds�Ĕ���U1���ڳ ���D�E����V`����)T�[\0W@����L���X���XLT�V���*��3�bV$=f��l�>�D�#���RTӪ�<;vaL��ȧ]*(��1��ZG�ZE��yL�:���g5�&'^!��IB��U�쉘Sx�\Ɇ��� Mp�T�Tg(mm2a+H/��rZ369�=���>=�ʼE�#�֓jp�>� ���5(�>d�5��9�f��etl��5�C��Q�m�WK�.��S�	��ACDv �Y��>���J��i%[�2���?��"�S����vO5)�{�n�z ��`ri�.s�b����I�Z�8���x�3O��5+�h^*���w�a�NRU�emO�i�{v������O��S���h'�2n&���o���Ȱ��`߳�6�k����	��oĨ�ץ?5.9���ș�����~��ۈ�ў�c/zD�H#fɵ;��� SmU�=m<�3f�V�
r�W���(�����~c���z��Y.��>^��?-xϦ�����S�)�wl�c��R���g�;;S��ZLt�y=��> ��3k`7���w�z��/��R�R�����`��j�U�@.�cV,ĉ��=�4����"�/�_H��JkW�unk�L�}��y��q?~|�F�$��Z]�usHe�*��ĄH)�4�9�3�mkA��	���T9��@o�lsO1RV�V�J��}�r^��Ο��h�G��f?^|��:��B�l߶�3��5�d{
C�*�~ե8~E�H9���(f�g������9`UV�mw<���V�k� S�Q���|t2��|v�Z�mOQΛ�#C���Ԧ��:1�1M��Ţ0��Ҏc�>4r��E&G1�B�����i�MY�B�9�2y�����D,҈d��B60�S#c��Kw}:�f�`�\MOI����O�Ё�Jû�Q�9��
P���t	����qʱs��hV��>��Su����(0UF���.���Dj˭*CI�2�f��L�mh���:u��b0]ŵ��NY{��p*c:�O_}x�a�~�Z���^��-G6%�����wv0X���ӓ3�hr�Lظ�����q��7�W��"�	cz������K`�O��~��_�׿��$
�<Zm�
�:V.�
0=�"����,a��p�g �I+�`���@�d�?�Xx��q|�s_�o��jkW��ex֯]�TR�#A����L�l!K`:gb�$b,��������a�Uj#L/��uL	�y4�ml��'l���y֙2�upp �EcJm��$fL ��[���_�%�ڵ[���_s�w�װ|�B5*2Ɣ��/���{�N�� ��E�ˊ��x�q1���t�`��7x�K�0u��?�i��"�q���c��U2�S9?�y��j�M��d�~7ݍ����GG�RB�9�mx�_�\F{���޺e�����ņe�RY�����,�7қ�[��H��\�&6��G6�q��/EfIEE����ZC��{(�
F�D������͓q�����%V�8�'��S��>!���=IZ����7Q�?���	9X�	L��E+I`�Qr3�7_��,p���hL�d�Vo"], ;W瘒ump�ۚv�$]�j�
YF��GM�1�k�Nf��lJ��dL�"�����3'N���S}l�jM�c�P��FQ�\���|;J�O�hr��ka�tbJ���)���dz�P~���SJ�{�c���3�����ً0f-ɈS_Q1�|���(0U��v�K��<�5�V�}��<�Hb��v��:z��[K2u:�;��mFqo�"�(K����+��T���w�ϒ�p��L�/�9H��{j&d���+6�X^P�~��jH�	+�z�V���2���n�2<�����~�_Q!��z��#r���;��k���I��#�|�ø���g�nL���/"��!�I#�'���o�@㤤��5�
0�T3'
���s��>� �?31�~� N�_V ��z���Ym?7����0�}�`#,5�n�j�
���8{����T��C޳�C�G�BP7bR@$�'0e�p�=9̩�8xW�ȯ��.%��gإ��_d(p��G�L�3?��o��&0UFX�	�?�8%
%�[�F�rY&ITg&Ѫ��a�(j8��#p�i���Kq��K�d~��\F�
��'ۤ�F��ƻ�a�}��=#(׺h"-ƈ-��,b	��bƹ�z��ݢ�2�.�׸/����ГB�)�3�� -Gѱ��s9,O�Ř��b&�.��╾��+�Y�c;M��������g�4�1E��dk
}�|��q�q�U�k�n]�u�����ߛLg�K�2��y~q㟰����l���Z�!!0�g��fQg^+$��Hw�I%�MƑ�+�L	��i�1e��M� gƧS���,�sV<{T�Si$M�թZ�v����4'��i����E��Y�(�-W@`�S2��\�AJgR"�Q]T,�HQ��SJ�����"�P��q,��p���)�� ӟ��(�x����̢�,pT�l���N�͒i1����*{^����RY�&�7�����a(]��?N>~Q�Z�q;�'��-ly`�8����kV"��zU�\B�Zǜ�9H&tR���L��K�*���'��k��[~�'tj]��w�aÑ��sp�	���f�"0�;\u�/�vbt��t�=�Y4Y	�ԐK�q��>|���`�c#b�{`>��y�YH'5�h��bz5KVY��>w�w����F����^�N��n���rd����:�w_�)<y��|�"�_d�.�zO���U�Ș�+h���_z>t�k���g�r�MM�05=�#�,v�_��F&ثgR�������|[���ŗ~7߼Qܸ�Y����5X}�r�cN������������?8�|�L
��I�O���C(�����8.z���*0���Ŏ�����O���D���FkǠ�o��Z�t=�
?�����'�x�B�=��x�9oD�����;(����+HbK�B��^��}�^��XPq�� b�As�ހ�hlW�;>���<%�֬�)��)����z�9��T�L4��}�'΃,�9/�#ע'>�jJ[	0C`:�o%���10.
�栙��W�N� Ɉ9�ԥ�Q�9=#-Jy��:2�>�� ����5�Q�����1$�mZM`*=�f^ r*PJw3)ċt�K	L6U^����Jf؏C�\AkrF�����v�����bG��ѷL��g��zb�$U�|G��l    IDAT��E��y�<O>���>� �5v��^�^0���
���h�XC�OP�>�eF�H} +؛z/�W�*�&ӵ�G�,:*��ޠo��I��o=)�a�t�j���G��y⬋�ȣ���������Z����0\d |�JJXp�9��s��#�)�*�6�i�D%Z��p5�Vg�|��N��:Gdtjh�&П�b�ы��=�8}=�2
M�4�j�-s M��3�gh�F3`��]���6�����dM�,�N��g�P.�^��2��=�d�˧�z��ֶ(sr)"k����FU�:� �������|�m��}��Z�V��>1Kuȏ���{�+IX����0���cc-l������y�T5�PZ/��o���>�*��պ���m�%�7�J��j�2n�0��Sg�>�3����=Ft;j�'`J
������r��ڔvZ
H�%aG���i'������~�Y ���dG���4�5z��?B�y`�J�d����k�.<��x�d���2�&���'�H��Xs�q������L�'�_S��-5�_�����y��f�20؊�?��v�-����|�����k�>,Y�lՊ�^��-�80%B3�Ds
�����x�)G���y���ٞr��az���%`�EAU������M���TW̏&f��w�e��[4�it9�.N�#�V��E2�%��1��#g�VIb������H��]��k�Ő�ŴǴ����X L�z��~yɗL�h�`�~y�r�|&�\")��-W����Ϡ8<$-S2�F�խ�Ԋ\��'��,gb;'ׁ�m"�qA�q1?�����c���Kyz�#���o��v�X�H&��æq`��kL��}J�"�p*���o��B�̄�i��o}�߰~�BaL�����������og�q^���	0�K�o�43�F��9s�"�J�U���d���Qצa4��!.�������q�w�]ic�P@"Vǆ+q��o�����T��g�O����;W^Jy��#�`��a��y�5+�̕x��=b���ĵF�{v�È�F���3	���-}������8��������'��iY�������}��Q\��9󤧖�ʪ�Q�d�Q��V��Vi?���O����KI��癘�	ZFmb7n,�'cb@`���G����>�������j9�s�q��rO�|�[�§��sl޲�fŁa�$�	��JC8��F�Cib%pɻ�"��Hw<���v�f9Zr�Dj�\n���Ϩ���`���[�/}?�(Cx߻ފs�y�nj_���K�`ZC�LH�BX�Ѿ_? �	Q�zsV/0=\鉑���.ǳ��}:>���h���X�|A��p4	�
�K3��jb�u�}�842�����9Z��)�T�k��YD�.6�tf�(fƦd]̛��E��Q�L��ڦL9��{+�+uaL[`J�4?w�b5��Y����C`�B���Č0��̓���
$��x]yu�E4J��T��r]:�ƪu4�&�h��/ڪ��L��j~ć�;0����C����GP�1����Y2�����$��{�F��&K�g��
�z~�~�v�N1��[���%H��9s'`�+���ēc]�+`O�DZق( ��������?� �q��'c��B�������6̷��H���}FZ�U��,���Ö��~��|��O�q��rf9U&�rsI,�6.U��,X������+��Ϩ�
j�c(�;X�h �|ѳp�I�c�9"}d ̬���
�N�
�Y���8n������-�7ZE��>q&�t9�b_:�B6�E������",��:b�Q6�^������D�y%�2+ӛ$ƞt{<tU ��&KEJ+O+��פ���P[����ٛvm��Iz��3�������ᰘ�s�4�?��B���X��Ad��������<S"�h|.,���S/|'	�X8��^���^���&�]bn��^&�DuM�ts�S8j�0�}�:<���pĂ��{��Vkr�q���娓�4�F&�����[q�wc��4Z��(�L�CS�d��,iaÈh��!a��@_����	��=X̝lT�B|��H$2[\��	N�D�z�Q�w�ֺZQ�y����Za���ֶ����|v��V>���ʨ�&b���f;������_v:�b��
�(0�=z����瀩������~�������ph
��'0U�މ#�������q/�ZTp�U��L*���V''��)��"� ��yJK�-}���c���h �E����8j4|l��nw�*�@��u���caL	L�4�T1qp������kH�^<9�\-�:��v���v0�u,�s���7ˈ�'�l��O]�w8��!����n��:�Zy1?��$��/���e��W�)	n�?�4��.cGu�Gη[2#�>=�ny��:���b����"�K�qv��c_�&�>��8�$�����ik�B?��;-4�	��|�]j�w�Ϻ�6��&&+1ʥӠ�p�ܻs_����Ձ)-��M�?�H\p�9ذ�u�u��i��/���e&��"idr4�u�7�
�3O���#�X�=�c'�>��siMD�)�*8���1�����?�7��s�u���\|�۰��%R�s`�q��=�80�Eah1�-�1ҋ`5.J��B���j̠9�o"0=���+��,|�oU,���[%��ۣ%�F'���>~����o|W��z��\��WΗ{�������4>񅟉+o�G��"G��\œJ�լa��>̌���8.}�?�U/X�%7v?��fx(a
3�Y��kF4�
ꡆ8�-������O_�;6mF:���'��[^�bVǞ�1ݼ��w\�)TbC�v�Ly�d����=r'���J�Z�M�<��SQ`���$�A#L�{�0�y&��~=����|y?=u�����K�Q\+� ?o>��d�C(ߗ�}��v���&��wp�\�������iYτJ�ذ��x�jw�֧gЮ֤"W�7$X��#^ȣ�j����L�&Z�%�3�є�K&<Wße�w_�l�dR��W�í�,�� ��	�,�h^��0g M��L��������#$pFc։��Tv��L�o�$ƾ�	�<C/ �?�S}C�ga���|e��_&@8p�d5: U6�`70�1Y��-M�̈́�׾��z�^����TXL0vP� H��<E�_M���0C�i<��~��p6P�[�۷�G
LC�%ݎ����B���k�)uo�)�I�)A�%��#)8!0՟U@��j��k���i�Q�"A�Z�������������9g���9}9��7,��>n�ź���=�ڐ��Ï�$�����|��=4�f7%*bIq.�hz,ds9$R	U�H���-Ђ����8�u��e��=�jR��ğUt���VȂ� Mօ�ws+-[;�w��
��@�0̔.�~>�
B �
�Dw���X� �S�����齵�|�LV�?�f{V㾭c�e�YQM^K�I��j�����,�DB{Y���Ѫ5� ڐ�Q��@S�h����:���,©�W���ƚUKp䒬Ql�μ �{LrH_����eǓ��έ��]�?ZB��E7�C�'�Fi$�������Ș�`��J-ȸ�5�~"���o��w�0�]�c���J����q;�����p`��B��L5у}��
�=�b�M��c�(�x)�<��]�
�i�x�K������1%v��:|�:���Ҕ��u.n7�cسw?��Fl��Q��`���L��:����r�SJyy/�Fx��7!0Mcʶ�(0����q1��6���4�������Q�����^R2�Y�"�Sf�bn&G�6�l:#}��R��Q��K��3���E�J�]Ot�BdD���B,Pp�;0mL`iW\��t�`0.h��,��>*���FV��8c��S`]\���>SM �n�c�|�q�][���Q�A}j�ʈ4C_��Ob��s`*s.ُ��7�e�N<�̓��?O_s4��I$8���ِDR�+�ҁ�r������O(If+�B1lyx_��z���M@���|�8������_��)���o݅�dF(��v�Hv��p�|�7a�����?�1����bhp�L�B^�zB��AW+�gx����f���������6�[����O8�8�s�� o�}�8���a�Xš#08w��m��	`*�"0��hԦ�.��_z*>rᛤr�l���Ƣ��c =H2���V<C`A`G���W}�~�:4�5�j9���+�r�p`V����|�s?Ɵ��v
��!q:f���7��c�1=�G����^���(Z/��KK���t*��R�����ZLlx�-�j� ��)C�w�n��'���6ng��;o}�Q���L`z��5��`J�4A`�4`�-�ޝȬ4�A�[������쨃��ȉ I��OE��GD�	�hR��L�)����{ԝ�L�l�I6&V��c
h��`�AXOđv`z`�dS)-����A�Sq���qɴ���"0e�2��2����
y��*0�yQ��j�xi�Zd�L��o�+a ���c�D�����ubL��>����9��Y8�r]V-�y|Q`���'� ���#`3dK��ы��z/�,��Tgv�����a+�ɦ'�׫�L�d��������� �SM�%����	��P�v���*{���BGᠴ0�!hUp9�z�nCU�SӠK��ޢ�8ʞ�f-g?� <��Hl��LeOu�X��z�U��P�=+�
ʹ\���M��<a��J[I��ˬ�<���x��u�sI<Y�C5�F���h�Է����g=/{�YXud?��ࣼ��u�ւ)��=��b� ��}��6cӽc�H����Hf�Hg�H$	T�2�O㹮�]���3��0S�hA��Q���s�Kig'�
�~�4��;YS�M5����OC1wD�j4e)Al�EhR�oE
9F�+K��"呩:�[�<q�=��,3+��?"E����~���n�;�ӫ�,�y$�<���sG#��oKb�uc��*"$��ˁ}?ؙ%2�.�&U���)Œv�"�ahՐKw�h~k�[�S7���c�����b�Lhh��;;�u�U,���{ݻ}nٴwo}��G��F�������N��n�-��d�T��ʝ��AG�ֵ%j!o�1�#w��㪤Qy����d?�y�y<E�0
{>(Ri��>ڀ9��hW�I�Qi�.�D���QIG#:���
��q<}�||����J����S�e�]_�s����x���ЮQ���w���O��d�zB�i��@<�>�i�L
�)K��UR!CL�T����b&��X�15`ڤ��Z/�Ԥ�K��q�Q>^��<>�Z�,��&'�ɘ"�͈��q�H`���#�J#O�]�`���3e�����%/b��e�U�/��b�ա�U��`cM	L�Ǵ>�e]|���I+'�#��(0������V^zL�\�<�4)0m5[VY��`^���
Ni<"���	o.ݛ:*�OB�6��t߻��8��a�H���]���e��:�=��<�����k���\�>e������Ђ6I�Z(w[�jѮ�d
�O��{���k���7܉X�+���T'�Y��N^�L+�6���)��/���LU�b~�^H�d��T���J��e}
��=�m�E�˗/��9s1�q�e����)]ZJ'�r�rY�~�X��_�x;�p�=��8��U8������-��{U�w�?�s/����꛳D��	�iT����G��f��/9�~����%(W1=9-*�Z��r��F��\.'�BtS�a�:"����G&ڸ���Ə~�kLON���׾�	,_�L2	c�X�~��-O��I��7�b_�zpQ�@W����(����A����#^����Wh��P��n����y�l�2�Ke��y�<����S��7�/����R�Mw=�O]�%l�|��y\|�����`z�N�O0��Xz�ȃ�9%�aM�̃,%�"g��S] 2����1��י?H�5*�q ����Sr�*L��V`�m*��?4�Śٵ�F���@. S?����	�ؘ��L���S������N�\��[�J��(0��P��Q� S6�G�R�F����>}_�n�DyV�&Z쁳��I%d�i7���:i2��6��UcH+tc�~C�\As|	�I�� J{��u����c�=b��!�?��ԁ�$��*"�Iѱ�D�V��D�~�G���,���=Z d��i�3jD�"
צK��%�m�=�����H��J�޿�d��Z���~�yƙ�����Y���?��޻ ���M����	�%j��>Wt6���8� m���gR�a-r������`� :���)�WäzV��)Z(V�2`��X�^��+���W�Вh��QC�QBy� ұ���9g��׾��8z�P ���+�J�/%�m`�<����[�����d��v7)&2)�O$h�B��tZ\��M&UmA?>S=���srY��;��L�m!��9[U+�O�Z���Ou֭>L��I�ƙp�j��y����ζ��pcף1�^��,{�d�����ɕ���Ѕ*O��2ě3��	gэ�6���E��[u�:F{�'�����d��;n+c�{T�)�(����g@Յ�&�@#�a�Y����=:�d���CE�l������5�g/t֍�2�!����Gy�4Uf�}��x�&�q�C���Pk'��(��!��H���0^ł2��L��R�S��E��o�7z����|�zLe�_\��?�_~�����kP��RV�G��YT��H*�@ϛh�wp�H+��/�Ԛ�e>���f;�X>��g?~1�^Z�\9��\9�C���瀩}:0-�c�������q)9S��Ti��$�\��6R	�(�}�c�N`�q1�?�*�MNI�3ow��D�sL���s�i^BƴH���`Z-Qʫ��|)+��2s}o	���A�4�\:#&J�J��Q���R^�L��ӸQ�M���Lb/y��u���4�ksT�V���߂�+��k`Zu)�͏��?�����H��Jw���V	�u���	����x.X��R!�;m��6K�@es�\�'�z٠,P�w�ڃ}�kx���8��'�/x� �y���ޒ	���A�xh��:Z�j�1�h���l��[A
�N[|�����tÝHT;*�M�q�	�q�o�)��������G����q7�*	dʘ֐Ntd�)k��%�y�YRP�tض}'>����6`ɒ#�h�"�579�({P$�j�&`�Voab���c5l�g�7.�'�?����z��;����;�L��{�L��T{3�w�����dL9��S=�׼`>z�ߊm��Y��6pϝwc��[�I�}C�%Z���Y�X(�` C�(�88�l� �*���|�q��q�w�Y��u���|K)`g�u`��+��][�D��B��0r��0��@�Y{1�扱C(��t��_�V���'�>��淾�m���0V�\���:J�(ͱ���f}�bd����9�"��G�ǝ���w��=l�
9|���wox�n�d���YW`F�w-�E�AGz���� u�~�$O����%O*��}h93���p�'b�`��
����1V���� ԃ�Ahx\�A�T�d]�8,	�f����̯�b��H>o��H�HRk`��(f&&��<�p��1e2��i��Q/��)�)2��S��`Jf�:0%��7�b����_������]���=�NIePXK
�ap[v���N!)�0!��0�c��Ig�4M��"26�-�V�-���z�D �=���'Qfnv*$�Ъ�Βx2�o��]O�5�5�D}涌zU��"q�����*_S9����F%�~�	x�f"з    IDAT�07�A(m^@���e��SR��܊B)o tm��Ϥm�g�
@h�`�w��v�	��v�X�N��Q`2�QE����vX�s��@i�}�<��Y�=y$\�P\8)��|�)���TΔ*Z�)T�GЮL`�QK��矅�mX�UG-�p��	I� ��o�/�����g���{���w�N�ص�<�S�6*���PJI�S�S�K�e�)���3@z�,�uE��S�_zer���$��K��/#f4d����(��(&P�� b˂���������R �te�0�!C�+R���D	�,��c�z|g�L�o�G䑋[1�Lg��E/c��8�	�cĨ�18蚔](QSD��D+���s�KCzG��j
��n"֮c�����<�/�q�,��'�ƱG.��y,�T�1�JQ�֔i�k�B�.����ݶ�ڍ�r[�V�"Z1�|�H�Ls�yRv���ar�gY[-,����\d�m-qΞ���"a�
�L+^�����H$�
%Qp����R
	���5g�����F��.yWECZ��~Y��m�!k\TVJJ�;t�5�YF�;���LW���"sL��{�
}�s *m�͗��l������4���>�ə6n��~ܲi'v=1�C�-T�I�jlyJ!�c���i����tse��>�A&��q1OL��6��|0�($�=AeB�͏
����c��̔���g�A�Xx7`J��xGp̸�eq�R�RSGQ�������c����C�)c$�K)̱wC�)��h���a�����R�S���`᧷<�/|��t���r�
#��D�^�d�12)3&�ZI^5�����"��h�i�4Tb~���_{9�Y�0���J`zɕ_Ǝ�����70}�q+��� �#���q.�u<J�J�:��L�[�P����j3�{�>����z���w!U�a���D��.���/<��#{]y'��}�:ܼ�	L�cHf2L[�:R�6����n).y�k�rqN�A��;v���� �}ͫ�l�R�Iє�H�`�W�VU�ll�0>]������
[�#�5����'g 1@ο�Wܔg�������dL���\�(;0�҈��6��cڭ«���T�)�>�au��_��x��8��(䳈˃�DF ��	��	����$MVqp��G���w7m���C����NZ��]�	,^��>Veķ�.ᣟ�!�޶�vBS�q���7�l����T�8.���^��uڟ`�����W��F���<�9X�b� SM84g��(A����ރ����!�L�PC
�mَ?m������>|�y��׿��n�Q�;.�$*qs�M�OӬ#4�Ҥ��ae��;�e�
�x�T����|$A��)��դAъ�N$ �d�*��_̄%�mR!q��T�)o!/��GLo5�A�H�cq٣�j��GP����o����cJW^���J��R��;�>"Jy�1�Cu2�U󣾢0�����F�v�zә2�-&�d"�c�C��1�eS2
�ܰJ5� S�;L��;1 SIz#�l?8����Y?�E��RZ���u�5`�5���`��Y5PI��}It}͹�lP�w0���[L��ɐY�DZ1A*~1�S*�s��s�԰F�dD�g�W7f�@�J~����p!���E]k0�S���ZcV=����>T�+�k	C��qp���AIBf��W�Yk��N�1\�w�&�w�g*�i�|��N���𿲺E��L"=��TOⰯ��S-�QTR�RgFq���t$D����Z�)�cu,������+^x6V��yH��%*Ԩ��G���L6�a$h����c�72�=�'��=���~�MUQo�yȢ�')#�>�d�WZ�V ��g3��=�{��\��	�]2����G�n+\�p�*����O�,L{P���֍e�,���M�<qq� 3��s�gt�3_��1�^c����d������N�n��{	=�3g�(wg�¯�]^����G��-tm�y�dNBy��"���]\v�oT���e�d�\�b1֭^�UG-Ɗ#�`����6Gf����W��C�ɣv��N��&�����>�{�=�m=�'LJ~�$�Qf<۳�KIig�0�BC��WL�����jW���W��.��M��%c�����^yB`jOӾ�l�?�I�?�Ί�����q&��J�������Ø˺s��!\{,ƨ��ݨ ٞ�Pr/{�z��PL�s��������Á�������������S�����b��q϶}����*1�1T(��%� 05�:���$ �e��c�@6�6���)uaL	껨�Z��s�]:�D��L�L��s�6*�S"�i-�\��~$��31���I`�J!ŸW�a����(���[C�8Ș}�ɘ
�x�v)���`J�#�9q\u�?��e��1�s�&V�v�=�R�;�-���Me�(���X�q/.d��T�ݒ>I^�11��Θ�#3�ڕqĪ#XXl��k>�c������?��򙫱s����S��睍g�[��o�M�'D&�"�h����F�%T8nDzն��=�`�w�u��x��w#ӈa �G.�ŉ���ކS7�T`Jv��������;��L�����eR]�1}����ݯŊ� ��z�I�w�}x�󞍁~N�_�TҪ�s���M,��#|����ß�$�5'�Z�K�;�G�4d�7n��[��84�����#�?�	]�4�3��G��3���Gd���*�Dib?��O162�W����?؇T&)=���)E��c����У���{q��mxh�T�5��]lX���ڕ�7���1��v���_�1�ڶW*��1��bl!	��m�1�c|�ʓ�D���ކW>w-�̸�8k�����t����`xh(�Z�f0:K����ڸ����y�Vܷ�1<�s7�?���i���K�Û_�b䤗U�MT���_�zr.��,��סg��#�4�9#����=9��ը	z/0%��M���ʨJ{��DC��8r�H{Km�e������a��he�g�*��ˣ&��ƢD�}:��4`:��JS�H��0UP�	���G񰊃�[2���Q��F��km��:٬�A���q�S�,nh $�]u坮�;ÃQGd�r��M\y�����5s����  _� �{S��S�C�w39U��-��kH��I��mր�������y9��_�2ݠ��' p�gmY��gV���*�,��G&e��H�Erj��`J��$_ҺԬ�l̏(D,����L�4񓂘����"�����On���������Nф�Vw�����5��S�Y컳
�Q�-����R��ʬ�:w?+�q���mD��c���{��>ZzTE�7�9H�������4:twVe�JRԹ�q�7�%��s4��:=�X�������Ex����Y���p�Q%y	�JxoVX;j��r뒡����ph���{Fp���p��[���j#�f'a3$پ�?���l��P�K�x2� X�U,XQQ�l�����x�t�Q�D��+��A�m�F�{�s��5�r"~��j*�q�~��[1J!�u-���Q��w(��"}��v0 �U��z����:�k����e�f3&޹n����\"��+	�7���5F�L�oi7���
z����n�k�;�h���a���9vN^�kW���E��ig���"������C9�
�r����u�}������L��%ifXD7�>R��)��:�iP(�lH�т�����B���Ϫ�0�=啥ңkQ����~��f9��77�جKpV��%_� '5΂��n���������RO��X[_�֋7�&�i�=��m�Q�H��mO`͑������W���3���"fd�̌�9Ѣ�S����_�1,d�9��mp>�-ƪ�Sh��hb��[7mǽ۞���'��@	S�*�:�Gwd�1E!��9�Վ��Ҕ���Ť�wj��������ΦPg�#�]����D�Dy�*"�D�\��g�Nf�L97�9;��,���5@*�Z�:����$�`����2V�Φ+�x��/ڱ���.�Լ�:�D)o��dsˇb�̿�k���?����:���H���&(u�^�j|�=)�.��^��g?���Θ�λ[�B{z��pݗ?�c���<v	�-[v�W}����s�>�~�sp��c0'�F\t��cI�E�x���hec��$�2*���rY4w޽�������i�Зɡ/�����}��{�v�J	x��z,��~�����M�c��@�P�E� +3�:%<���q�?����z�
������f�q��0o�l~�QU%I�Tg�r!H��%Pi���o�
�����dX}�<|�����ʽ��ɂ��[��K?�љ$���(� qv�j�����X�Ӽ�+Î���V����QS��"0���m7�*3A�~�3��f8��i6�ۚ�1Yi����ɍ���{���$�8u����՟���i�ʏ�>:�+��s���>4�id�}2�	o� �<�&&Ș���b��\��Y����DڈQ������k֮�QG��~��pB:���h!���ul~�Q��;q�-����'�춰`(��.y/��e�@�������I\p��QK���SG����Z�F��ͰcD�G�`�>0�0�DXO�ʧs^���)���U��@��������aiU[��3���̽?Ug׼�ɫ�h��2}}��*��NU-Xb��?wkuL�?$R^&�Cc��T�ܨ�4���F��)tkM��U�7��d���q1��K3&q���k�l6�z��������I�L��:rY�����$% �:�>�&)���qeLSf�入 14��e{ҧF`j]fȳDB���'�nx;#hęJMz�RY!���E�ȿ��#�?�i��L�����s�沊�a��SO�������B�/#�%��eyR�j����y?µ-����ߞ=f��'��C0��b��T�I4Q��h:�sG�^�:d���&?#�y!�Ѣ	����V[�~

:�}%+W�Bw���� AY��/-���� h�x���
�ud�$9�I@b�k0&�b���ZG�2�Nm��8М�������pƩ�p����t�0�9 ��exԘ�� -'����{��8p��p�-wឭ;��QL�j�Ē¤R�cKO"�L6'����:�5��%!`��I���q(�'s��2�f����:�H�톻�@Dg"}��s��|� �ݏ�:J�j�������L]�_�}���Z�����,�K�l6gc^|�Dzn��JD�<�����)�1W@j�����$�M�[-ԙw0g�� #" �n��1����Kb�!�bN?e֭=K�З��e�C0��a4��UF�}˻�ǎ�����>�$��8��~$2}H����CE�2�;Q��b�D��F�y��u=���33��X�������|ݓ�=�Q������zGx��xгǟ�j�%TE����V�����d��(P�~�f=W�V�VK���\7	�t���LaN������u/?9�Զv�s�Y�G����-����Su��a+�a9�]e&i��my`/~q��{�&��L[��J�+�]*5)�RN0H�ev�8��*�K���xKƔSjM!�K�(�E�4�~|b,1�P�O����Ea���4�doinpP�㑰b_�%-���̒p�Ou��0qse�$ �t���ncK��-�J㚢�����4�J6&�b8��|��8����H���S��X�ӟܢ����ʫ�.�����|2:����iq��
Q;�V�zY�ik�I,���c8ja�,Nv[7ݳ�r�q`|/~��x�+^����?M�.K�dcHSf옰/�FeV�xX�bJv3�@#��d�x�|�?ă�7)o����v	��ũ���1`����~�ߵW��3�奿��T�%sL�s�q8��_�%s�&����q\�����>+��٣���h��j5d����d2�G�\�t�8��;1|�7��_�N��Y6�\��8y�R!�!׌'p�=���߾�љ��ad�}jZe{�Pd��bΕ��]ڋ�y.��2�6!r�Z�f���/��g4�3����'^�Ճm�������~�;��׷�݊!�i�����/�iIq#l{d�������H0U��m�SIqޛ�Ce� �����L9��_���ҥK�?�op� ��; �͓��e�'��U��ֻ��_�l߅z����y|��s�k��&#����৾�fjjݜ��]y�:,U"&�&#�1�F���:�4Ɲ���A�]	�1:���SV7�0�e�[9^7�R��'��`�����}��A��R;���$�f���1���V1�VhQW��/��ʲ���7�ʩ�:H�&�1��c��a�03�כ�&<�y��3���f3&؀`#L���$���V�suuUݪ�=������έ��x�����U��s���������J%i�E�T��E��ZAcע�1`j�*�ɘ�J~(2�� v#�:.�'�)�f��^�ȈiXD�t��d����4�`�C��Q��Q���T�B-��n�N��i2¨�C�I�S�8���S�*�3��07HgU��x�:������LmdU���WU��xҤ���t$$v
�^���1Y�[,t�2�`����Ӣ@t�ǏY���J�|�/gj����:cLw �p������k
\2lo��aZ�O�,��?K�,�*���r+ L���P�	`���P��PV���Ǔgi�:O�umi�	ɪ�4��ڡ�W����f�c��.��a�>��(�Yu�5i�9�jo*ea���"�W�^#��a�9f�o��jb�Q/�pٮY|�sn��WµG��K$t���T뢉�'��h���^3A:��<���<�'�����x���8y[���b�a&REڂ��T�`��6�Z�j%�������s��d�L��h�ky�n�%Ru�{r�S���$T�Zr}�Z�6Ռ�*�B����1�	�I5�?�Vz�	xEN������1	��Af>(��{Y�G)l���x�FF	B�~d#u���"�'2��g�W�z5���i�۳����p���8t�.\~`�����J�i���FUM&:��#�N�n;�Z��w܇/��x��h��(�fP�La}�:�h2���0�ehf
��<��;a� 5�o���B��M�)$����T�����0U�W����^ �͝1��}}�4�e��.��?��ns���W��REA�A!��B^y�l����=颚�0U��e�=�_}���� ٳM��I��甃�g����YP��y)�Ͼ��*�TQ����1>��o��{���ծ�����N4Bo0��!(�Wk�cZ�c3��B��kU���7�)�)�>�S(�M#.���%7�Z�h0Y�a�Tr����FD% il]��Q��W^Q��d4u��=��TB�P`����nsK���s�0����Xگ� 5EY[f�IJQ��c8`Z�6qpx���<��W��駿�$������QM{Lɂ�[�f�	���JӴ�cXb�C�YE��K]$�u�{k8���G��vX���XN�����0����bs?�C��O��q`iU�[�I-(f�k�D��t� ��HH����r���?���ATF%�ZX��T	7\���?�g]�KӜJy�=�����).>�d0 =E��>��a��_|�5��x�'��w�6��ۃ�va�^�0�#��r&�"�)J/�p�Ã��޽�񶷽�+��:>�Ż�w~ɨ�=K3���Y��y��WGd����/���o�Q�YF�^��<<=���Cƴ�g%��a�<�����_���	0�̖�q0�X��Uڡ[Q�Y㩭-�C�Qı�6>�W����GD��~����w`�v���.~�}�o?Bƴ*�W8.�����Z��� B���a��R#�������ɶ�g��Q,..baa>|Q�Pi�����	�+�x    IDATUw��}�/�3_�_����Ob��,��_��x��nA%L��kg�����q]˗�Ru�D��Wb�#����,�<��Q..}�iǇ�x��+a��;B�,@��"W�3�ZI�J{D�a4w�.�v��qSK��M��]�s@ev���k���*�hl$p����"l�����M��ө�K��+��L�1mQfj��$c��h"����q1�؆Iyi^Dp��a�\��֖�	�[�c*��� �����P6��q1L�)q�#>����*0����
����X����<��#��)�m�<*WդO�?ԀB�y!���d���#L��K��)æ��ƀ�NqiX���V�]��&T)�if,�n�*I�����A��cS���tg%{"��ԓV%���z��Y }7�=)���M0�i: k�`�s���t& '}��bA`��D���$���Ǵ��+�]Z�;b�9���s��N����d�����x�Uu�[��`8����ѕ�1#ʑM����Q��q��OM�m�6
8�g7\}/��F�r�XY*��,���iq�R2�IYw�d$<Ȕ���� 'N����8uj����s�pq7��͂Y/��%�i�TF���nfQ�ꊒ�j�a��"J�g^��R��Z����f�
8�d+��� rә�L�d�h����{�\*�V���_�W�J���Ϫ4O֓l����#爍�3'-(8�P���Fˍ$Gq�ʵ@�����ʹ�<���2���@抒��Ժ�*槱<?����Ɓ��8x�.>��Wf1?��E,ܗ��P�>d������i�����`4��v8z�|�=~O�Y��-��cJ���,�29��V JI��(�O�@l4���������}cZ���٧�2�oo����*f5^iϸQyj�Ɛ^8�X��~BODưo�g��g�C�����9��{e���S>�n �m�W�'u�eaB�><��H}���>��k��[߄�|�����{x|�N�P,���LL�����o�z&Ao��u�(ɦ��aEɖ~�ￊ�8���f��*z�1��;0b��ZE�^n"��:떤��L���������a(���T9aLu��Hy�(R��F����Z]a<�$a��Ř
���(T)UO�������P)�d,^��h��t~V�^�/��h)N�41*Y
��'J̡��=��r`x����������1���U�eT`�G]��1�	L��T彩\A%�Zy#�7P`ZI�����x;������o����?�fs?�o�O��X�*ɨO�$0g*���)#&QCL������ ��C���=�B�Ǯ�]��p�����_�Y�|��K����S����hv�(S��y?l���pٮ:~��ވ�ܸO佣��s_�G����:XY�=���cj��F��U�B	Q4��Zߺ�Q��J��_�5,-����c��w�o靡F���{%~���Ҝp^�_~����O������*51�Q�;=�(��Q*pXz����]�o��_��*ڳ�z��Q���)��N+�ل��גa����s�C|�S��?��� ,�������%��נfֿ��w}g�����'�1�WEjE)���d�L�^�^O$ Ť���7��_�Ί5��Vw�q;��ٍ+�<����4��H+d�_�!��\�	p�}'��?�;�����wq?�����"3�k�F����1����qeq��}n��bK%9��M&��>�-Oc��,6h��S(���E�,\���f)���eY�n:�����O:8�Ԡ#\Ŭ����2O4b�Cz'�:� bv�EM&D}���"��]^`�R^9�ݴ#Gi%�d<���M���m0 *e�1e�E�#�H\�l5�g{�q ��9�Q�;"=�L"���1.S]�0c��Q�)�#0-0�6�����$&�7O6S��?Jg2�i���dWm Җ�(X�q6���fP
���>g�S�a�=�yߩ,��f���++�ɒlk9�k�[����-][��<Z���2��.5v�����33w^?��kFZ~Irc���3OU�g��L:'��SQ],��Rf#`���rh3*��Kic�wgb���vM�m�9S)K�ȱ������Y��5��w���W�!����-�g�|t�wF��j6���
K���.��~l뉺[:��(�"�Y�ƍ�^�����p�Շ1S/
�jf���1����KC�i�k�J
�0� ]��C��M��'X���w���1=vg�]D?�Ӊя�3+�I�XIg�n�(�턣ު�U��(Q�G�EJ�eeo���<�|�PNs���	��Z,�y�^Xq��ZB|���K�01�Fe� ��
Rxa�Z�+�����!˕�+/����q-I����&6��&E�w��C�S�"�p��}���øꪃ8x`�����g���`�`)C�eDR��9�Z��B��P71"C��=���gp��������z���x�Be
�jɨ����;�Jo����43'�������~O���X�4f��W��\	�GCH_=���}��IWC\3(�Ko2�Q>��!�z�������|h�u�{�s|�x���yZ`*7�ܟ)�M���q�qs�-�������=���zmݼ#�j�`�vF�����%�M�^�_���K߇�,��8���l��_�w��֚C�⒰��>䐉&�8��1�j��2נ�-�B%��(2̓r(svz"�%0��D��))��5(�%c*�vF�N��L��4/"c��t��b�i~�S��͠�r�r	�b�~���:��3�i�P��Š��)-�K�- '"��!G��JB�09OL����q����~	��-w�)�����	��c�Ņq�|�\A%z�gk���|V����R���jT:.ƥ�ø�ܠ�ڸ�ڨ�����-׮h4�N|�������JP�����u?��z�4�&��(����W+�v������?܎��3x�ѓ���ػ{�jy\q�4��so�n�Lg��|����������3hv����d�x�-����ܛ����.�;��zW�`n�����9��y�T
덊BL.���8s~��{���6~��o�-Ϲ�*#|���x�}k�dY���+�醫p���87'��w>��<N�2��Ya����I�J#vVR[��xВf䛯ޏC�gphϒ�V\<
�v��?�Z�,�O21v���:e� l����}G�W�E|���c4�q	Ǹ��x�-7���]����������N	�8ΕL�L'K�E?�#G��>ƃ.F���7��/��&�Ct[[8{���.<�Y��'~��XZ���_�$�H�U��Ñ��6���l�ӟ������p��^��k_���u|�ᓟ�_��q�<��2����j���V'�C�A�M����e�=�����ٯM�uK�vJ6C�u��{+;w1[�T�Y}�	_j������J�Jy5P�a�UV��T�Ikͭ3�h0�3W�>���z�t���SVR)�ƴ�UF�ĨRB}eQz/�'}�A:��a�7.�%cJ�8��!�)A5�u�Ā�]~�o�H���@��I�fK��u����q��5y!yf<t�]IB2�/�|�\�PZIF�|��N�ETj�� ��f�`�b�8�������򖙨�^`�dm�(@ף�h�T4��fZ��3"_Kv�J%)Ҥy������vV�3�۶��%e;_/��)A4�JYgM���;d�a1�i6�P��o��vńgm����d5�	��8������4�T��$S�K��{*@�c���n�"��Y��K�sPr��7|t�nc��^ڝ�$�j��I�Y�%X�:w�=�Ge��A��q�A��OW�a��+p�՗�Ё�ؿo���p��{n��k�e�L�l�cRn�B)��pq8svO}
=|O�8��Vۭ�����=aC: �E؏ܘL)�0J&�[���P��.�Ĉ�N��ZE��Bw�\�?�"��L"r�vku�x|�>U)�RAA���x�x@3��M�t�)��m�9��L�[+�,���jL��Ni\[d�U4F����,-�a��e\y� ��� ܋=��� ~/�b���������ة��n	kŖ�g6�x�6���O��S�p׷����V����\��bu��6�1H�G���9���rB��G�p���p����f#���.�|ol����}���5�ggmq:'W�g�/�s]S�����Jl
s�U.�,���l!��[fu�K�j$��@��E�H���$tc�s�V�%�U�_17@q�Be���o�����EU�i����l�Ό��"�%��u��9S�y�oN�ݟ5�C�ϾI�{�]���閬�vD^�+�4�������U�1�	z!^%�YϜ�z�uu
�h���C�be��Q���$i5�s���|N��t���V틛2��q|�0�6�#�Xt�5���ʥ��y�n_���[��k5�1-��1��d����G�k��.-_��j��#�IT���rL��S��)���%�~�6��ӄ�<n��Xt���t��X1)�bb�.-���ٙKa�A��(B)icԽ��x����?�j4�Ҋ�Gy���+_��3��_�O���|��6�e[Niҽ�z�ͭ�y-��0����+��'o���MT��߳�\���^���e/}.v��$0>~��?��_����mՠI
��PeN�a�A.ꠜ���G�E���q���\o��?�7��嘝�˛�z0�-�|y����C��m_���b��e����"��ͻ���܍&&�E��H�V��S���0�A��Q�������LH�q!���#���rq��]Q�緅Q��⸇}�g�?�#��97aj�.We���hi���2Np��>��;qǷƅ�a;�gfE�ӏ���8�T� J���;*̠Pn�,W��̓�39Dy$�H����M"o#?��p��o���*9�������`v�&��r�+�	��^�^��N�6m�G%�5�����q�'�iu�b��<���i	� ��Б T��W��=T��ZC�]j���8=4Ryc`6,�R��$M�W������A�̖CIZ����K�nl�DE������~] ���6R�+��UJ�V��Y��N���sho4%)���q1��X(a��y�X���͗@p�)/]��V70��z��yaL)m��s�8�aI��(G*��ES�&��~~n
�RQ\�Թ�G5��n��8/l܉�p\�P{L����G�A�i�!`�{�I�����l��V�R���kR/q�B@��8�zL�����<c9ش(��W�5��q6��Tc3#4�̨��g�0Mޫ,�����=̦��R���O����98�ľ��+�*�R����{���Kj�z��]ā�������!cW&��]�qn� �n�ｩ��o5�񌕹�W�݄J������ܒ�	`���ޔP�����F� ��SUR��nv�hO���f�D�|n'��a�h�:��5�<IfT�b�ó�@uq>�����j%��v����W_. 芃���P�$� B?��i�5x��d�K *���8�xh��onc����v�ֱ��ƅ�[8}�N�\��Z�6�G�Ӫ�G��-G��\f���V�o-
P͕8�Τ��O����i߯���*�J���u�r�h-��x�qd�����E���T�4C)bz��C�biq�ru��+ ��,.�bii{�-cyq��U�����Z���5����+g��a�Wv�淚�3�]=~w�� ���oau�����Q�"�(g��*d�F:Ô(�/��J溋L�̿l���T!
x�C�{FV��t����f
9����a� ��O瘚ov�jW|�Bu�t5h!�+ʺ�Y���3;�����!T������>�ŕP(��(�F��Ll����2�X{4�����Q�Eh��V�y!�͏�
+��*Z<�*��by����|H��&_��
z;������1w�y�I|����&N�kc�3�1C�}���}�xC�)�	Lke1.�h��SU��-ke�|�x�I`ʢ�i�^�x����[e"ݘ�G�%4�@�� f����F(V+�zUW^S��}^-���BE7���"����Z2?���q1:.KH +4J�*��{L�=��tT����zq`L��[���ȷ��W.����/<���q>��_l���P�P�T@(��~R.#�Q6p�4R�P��LAn\
�A�a�k���C�.P��p���[w܁�v������ί��?�=�bi���D�7�l%� I�,��������O݆���B�WVP��P��Ш籰P���j����.l���M ��hL7?�SC!8�`����q����Ѱ����}K�ϻ�j�,Ncm�Z-V,�X]��ť%��:�٧?�}�/Q�-bfnj��^���VO�(����f}ʋ�|>yi�N�Y��M~R�dJ�̟�aʼ7tM��J�3`���EM,4�x��7��+.��(�W��x")I p2��d�ᩳ��sX]� �0P�5���$	{Zx2�+V1�UĄH�#�H���J���u&8z�9�5�Wy2>�H�u�ci���/߃=+3��������s����D�#���+hGclwbln����Ke��4�P�!�к��ҽ�fUҫ�����Н`����,��P2.%��zo��d�דv�:z�|Z�M���>e>v��$�6��>&2��3�L�2pc���ِOW\��D����̘`�i{�)�bfVQ[��q	�+��𓳘P�Q28��h	LiE�1��+���S6�;S+`��}2��6R�ْY�dP�X�?�5�ҽZs�Q�����M+мO��\t�e��p�#Me��ٹ�&�t�5�4e�kp�g`��!@��a=3 A��F+[(��b̮
(-�t_��W��y���Yy/��W��#���:��/]j���9`��N$y���yH�v���<|��}`,e��f:a�%�X�=�pz���������]Ni]�<����R m未�3�O"���`�~o���zR`�e_Ē߀������^����~>�?�����֙X�����MO,Y�+�d\���aV��`��Y���N����E8����d_�ʤ&���gٗBow�����c�NU�׼����E����`y���9�������"�4���Υ�>��?�����������>���Ml��^���zQ��9�k����3[u:��[-l�;r�t��!jc)�
�*6Ƕw����{�����-^����m[��*�z��2�2�fj���c����j���g�L�R�\�Z-ɿ��O��������Z)���j���U~��Q�&ĵ^j�A�����\��T�sF#��C�8y�>~�N�����]h���M$l�`Q;�FC�R��Q@�Y�%����[hF���k��\���B�K��^ �`"3��ρi��PT��
��tֺ-FYO��a=��v��s=m�H瘦�ӎ���h��A�f��m�/��ћ�p
ִ��M�����-c����_k�&�OD%�Ey����?���ś��K0EOI��jL�uc���;X���Lz`j�+e��A^.���|��������� ��Cl��ֳ@���\�L��瘲Ǵ"3H����K���S/�s�s(�:]�d+قD�E�m`z
I�(�)����,(坫U�{%nnk�)��c3?�9����Ѡ��u�\!�F��Ϸ�Rx��*:Ǵ8ư���T��Ex���GK�3*b��TT�q�zL�x�IyC_�3<����g�=�?����6����c�>J�s�x}�Qʎ�V�e5���zEm���U��9<��J~��h�jn�Z>�sO����p͑�x�;ߎ������t���?hR�Ő6� Y��\Nd�'׆���n��?�9��1*�:���1;7��8F��0�c���e���!�*(�k)C!M���R�2����.�Incؿ�ûx��|ϭ��ч������0�kkM,-����n��_�J|�ۏ��?���
�q�g�
<�,�|R�^<9�    IDAT�2{_X1��֌.�īj��f�~�G������賈B��d���p�A,q���4������2`��T���%2�����p��P�4�/���Ğ~���|�cg��&�̴![*��c"�K0I,��q2��v9ǊLs5���y�x�,̔1跤*O�����Eb��Opz��Sk\��K<�=EY���3�V٘�zJK�*{���������(�VM"�G"���J�l��-�}4.�M^e%���,���&����l��K�7����t��'���5R����*�i�Q���2�b�`2_qnVW\��LR���Σ��`:�� ��=b ���g��!cH�(����-��mI�X0(6jA�+�G�����T!��RY0RW��Ɩ�2`jc0eNX+��0#����Q�_s��C[��\=2�m�8'��g�n�a�S�zh���f�4���!�<q
������̰�ʰ���U���hk�FG��d�.f"�Z�ZIב�yZ��>�QU������T�&��Y̲�������w�Y�L�Wv7�k���V`� IF	�2OJN:@���l�KO��B�~�\����ŀ,
�)#[��i�ix��a�[�j����/�p��8b�T~,�i� �	[�����7��>T9C*���dl��zr���Y�Vl�d@W�<zvj��+��Q�<�Ԍ}�<�oh+
G��q��u�Zb�2]/b���ޏ�:�k��s3S��ի��+}��A�,�0_��۹���؝���@���c��z9Ò�5Cp���0��~<`����s��x��	\Xkb}c�� �~$��k4N(}d�'�l��>+a+�,LW`)���W˘�k`iqFڇ�.�^���L�j	�z^��(��$:�In����Q���Zc}��Ɨ�BJ���"�U��JA?c>�~46��h��8s~�}
���}8���v_ =(��)r?�Q�(E`R�tD�٭�"ѕ®�B��7�Q��!���ڣ�ݗ���9�����S�"�q)��KT���RZh�k��J��@)�#ty�1��H������y<6��Ξ��W�̰��Х�J���>��s�y�  ;BQZ�4�`q�� /@пK�&�"�nc��m���W�,�:(=��<Dy\��E�F�K�r)0uPj��L˕+T�u�ǎ�Ꮋ����z3��V�Vg�n�?,ɋ�`2�dN��2
��Jy+%q��`�=�R���T�K�c�3�����oE�j!��j�\q����D]�㼴I�*%T��P�UM����H�D �C`��DธVKs�jES�q\�0��"�y9��%�ه.�Cdɇ1����?;��}����Z ���w���V�*�Ҕ����׋x��q����ʈ� �5��K���^���@_4r
2��&{G��sx����gp���������x���<���K7l�������Ǣ���h���u�>z>��ϡ�JP,T����F�������*���F�6Z�j�Ň�@'��L$7�0��=8�d��������1��{n�ٓ�q�w"�b�={K++8ph?�祯�]����O��Ertql��J:����ʱ��KA��X@Ak��U+uT�a�֫�!"e!G��tQPE�6qh��u��ؽ2Ǖ�]B���؃G�cQ6��O��?�f+IC�TC��q3��ғO� ���C4Aт�&n(��#��lT���f�V��-L�\�Ͻ�J,L������85�"�����t����'���d� �>K�\S��ٷ<�j��~C�mh�0���F<	�Yɒo<c��������Y)8e�{b'0�Pm��^]�;�hO��J�&ǖ�d�li�������U#��ol���yQ��ĥ�%Ns�r�Dl�<�����ȾK���|��4��7?���-��-��0��S��cI��QZ)}�C���){L)�[s9�u'D|��*���:ǔm�i��Z���ǔU�/�Q����:󪴲qf !=��8�� 0�u�?!L���ln�'�´e��Ҟ�L$XVIv6�M���ED�Nkc>R�px�M�m����'�a|��>Ճ@��H;��������Y���L�A�|>_�V�wP+��i���V�}���DԋGA�i������g3&*�~{��)��9�g@�8���]w-)�d/��J&��B4�5$'	���qJ�eY�����Yb _-^���I+��I��=�/qy�.='��Y��#����EY�֓&���iā�:�� ���<�ø[żB����ha(L*��y��2;���O�S5�ݽ�k��Gđ+�#0�P��p�<o7ӓ���S}���O��f��%mؑ!�O&]�R(��9����S�1B4b�)��1�ϼ'ʞ��KH]nH`�O(m����JU<��Zi�G ��(�)g�3Ǎ�|NF)�!����iA�Y��S�xfrq'p�h"(on���las���f��N�Y�S���'����mD	M7����ؓ[C��=�°J�Q��� `3�bDU�:Nk���^<SՊ�a�h��m��8+w�܏.	�JO�}^t
qC
K����%;e]�dc�d��U�<pI���f۝�^v���>ML��Rva�X�;5I��7���r���+@V٫��d?9-<�\BZ�-�l��N��0�9�������qp��_y����b���Zew�+2��Sؗ�g���>�w'���O]�̩���v���>z
w�w�[�Z3Fs{��v��&TlQYZ3�0n�=�Б1��E�+�F����z��b�B^���6���1��-4��LC΋
L=��q�l�"�i�nc�����U���}�Jz�Ơ�J��,n�8�S���m��T���")�u�i�9�Ɯ��hb:���P}`�6�4��)�����.�F6��O��>��g����%���ց��K��m��8`٘T�7�ݒ�-�dz
4�ႤtG$>� �5�����PE���� �&n�j��=��g�x�z��p),� ?��/ɏI�xӍ]������<>���ͭ>J�����V��F_M�4�e�(0����Ԃ�e��s�W(�!�K�eH��9hbؽ�C�kx�Ͻ	�|��� =}�4.�m�k_�S��W_{����ã'���w}��vP�كh��{9��#�I[z��1�"�(I/5?���i\P��!�g�g�` �����T��<�R-�[i0ݵ<K�ZI�}1k��4H5)/���?��<t[��|Y*��rEzh�B� s�ţ,W~�L�-1�k`B�ɼZ�k/���^�纡[�����-��5�-��7_��i���W�5��G����y�@3�·��'N��1�Lm	��u;+�Є��^�����3cQ���4��<]M/�J����K�}����<oB���.iR���ġk{Q0;��X����L
�=��uOs��:c��L�~_p��$�����籽�!����e�W�T�˾sa[l��vQ�±1<�D�r��Z���0��"tC�.4�H�)�bo�xs�VOzB�WЙ�"�%8�UP��Ƙ�y�q�:~�̃� s�5wO�+=��L�-xL���u|���ʯ�<Iۤ��ȓ�Lk���	�t'3�e\�f,�hu^uv�l-pڍ�5��L�!ۿR�3�0�0�(��ʥ]<��:59S���)�ݹ���?Hqw����~B��^��oy�![�1����Z��3O);��#ui��J<�"�>w�<�o�u�U�T}�lA�{cW�r}D�cČ��W�\��*q3�R��2�^�6VC?bF�R��3&����ORi����Dlb�\@�d�n
������kS��א��~6��P�7o4����Dڳ���3Cf���ڈ�1W*Ƙ��b��\�ؿw������w�,j4Τ45ﮰZ����AKM_=mN+���t�������9��|؎�K�.;뇮����d;m�����&��?<^�sIcU��R��
5V8����&V�p&�����y�wp׷�'�`s����R��lm(I1�P�i�o���<����3�rI��)_ڈ)~H>c�#uq��k�f6�45�|����V��|�s�e�z6Z�(��Fd|i�sp�uh�b����aǇzL����ݽ߭"$^��^L��N�5�`Q��"��S`�9��)q�3�m�	�� %q.��t��o��-7�KKV��Ǒ�S�W?�Z��9��`K����p)0���ү?��W�b�;VD�,�>p�O����C���ٵ.:�<��*II7�Z�Ґ�tLB�\),*�_	c*�n��H=�:e�Q2�3H�%��T�i�����]�xI�t�\���ֶ�!����}Ĝ�R�֫"]yw S��e���u\L��-뚣j�s3�K9�8B2g�H�M��縘<A)� �R`��>6t���A����ݸ���?��]�����tP�6�KW�lf�Dt���S��J����K��!�8r�Q[� ��h�F1�Fa���9{�.�m�x�^�7\@�6������T�`fM�`4e;[E������e�7���kX^ڃz}Jz�D�H�MWY^��:�Ť�f��^Cn~NM��ym�0r������О*��T�d��%c����o܅�<� _q ��|+V�9���}GO�Pn,KPϓud �*��#�!�.�*�0�Er%>���eE��꼧}AtE졜�Qa:m����|��Z��t2�\+�Z�U�]n�N�G�8��<����b�(/�T�Kɱ0&�ф��dI
 *`T#��,h��f�Ze]Z���Sa8@i<�ũ"�;�/y޳�4_��eS�=DǠ�X���|��3-|��Gp�cO!��dLc�"���H�e͛�+�L.�W�+�A�"��tʔf�;R�Q��e�2�M���Bҿe����+Dk�~.(#��B
7SуH��$�5H�s�,��0�l-�|~��vH�[�(�帘U4�.�\�bn�� S��ׁ���
c�g6H��(�jc���R}e�麀��S)*��g�����b�C3?"���������0�UQ���9�L�ǔJ
�]Q�R���V��*��\�6WГ	�/I2��Y/�Iv�4#CKd� �!�w�h�M�O��3��T"���;�bg�3*�P<Чo̚=�����c-�$)H2�sI�� ��jo��^�x�K���>��Ui�/�5��E;T����J)i��s�z�%���f�f���S�)|�ϧ n�Q����z7%4�qY����r~��r�a�?�l~��mv.�]���)�nt/eȋ�L�
�����8����kT��� ή����M�B�M��A{�r�>F�/i�ϴ��ʉUf�\z��޼��20��j�*�G�$q$r�$�:����qҗ�����˳ؿ{I�Ͼ�Z<�k�����[�v#5ʌ�v&t���9�*��6}��=m-['���z��~��~�x?�n�ں����pn8ȴ�����L�$ԁ�T �UE��^l��x��l|��y�9��G;���M�#��i�X��֘#x؟W�5�|% b�
x���MA��+V(w�b�F~�������T�H\5���K����5W���R?H�f_�~?g\�u�]s��ٞ��
���rKO�Y�b�T��vIug~���Ӻ�_+�+��!�wi䞈�Cxk�W74�*���|�~OAi�=L5�{�Z�d�8��F�����mL�b�](�?�z��GP�}�	����j�3o�̿<��kF%����'�������8w��v?�v/�AB⢀�C����Cft̑��Ɣ-��UN���4���|U�ص�:Ǵ?�\���4G�Ԁ�S� �E1f��rqI$�_Q��V�:.Ǝ09��[$��@H"�r��:�n�g,MOӑS+~
�2#㵰�j~$���9�#�6���V�����Li~�O}���=X7��WB�8�X�U��Y�yUV�ut��b�~#g-��! ���dl�`�D�:n�*�o$�������F!j�k�����jo�ݹ&'!}	�#$r����{.�3�{?�Y��g����>��w�C�1���,L��]	.⺨���L��针�A�TļA푥b��F���8����/�z����=�yv���m�aai��Fy� ~������P[)����:�w�Li���2�\Dtn��@����-�#j5��So�,2a#yY1�Z5@-#�ph�n��Z�AJ�1�R�E�P��V'����ѧ���F;A�:-UO�V����3�DIm�UDEƌ${.��l�8����'H�:*�#�Ǳ4V�����xѭ7a�Q�d$�zrt�]�)�+�&˛��6���q<p��qQRD!�9t��Q�1-��0� -�A�oTC�<�Ҍ�q@6iD�\:8	��ʔ��p��i\
DvlZ?�����q9�i[*��X�=�5K�5֛��%�^�忩ѕ�
=p�|$��:[�4�P`*.�
J����>Oޯ~��kh^X��s++�--".�¨��@����J��fK�F��������Gf��`IY�9s��nwe���m��F�3��1�#c���R��oݸ��գ1*# ��0����{f&��,%�z&`j�V�	��,��Jg6}�L:-�RPO|R���m�DL�f����j��1���kL]��$y5`��k)�H�.��dC@������lja	��_�Nm�6���?�=)�܀�>M�U1�uj���?�O��m�By!c\ei���ܼW>��"����K�S.�aӂ�PG�(���a�������YM�����g�R��-7��RF��PU��C��'�k["-�y�S��4a�.;�VHuV��3_st�����w�ɾ[���Q$�:�3D"��]���A�è.`�]qh�s�8x�n�߷Ӎ
��(w굲|m��DnR��@<�i'�$�)�|�gm_��{���"���Lw��&Q�&�(S;��NL��<�,k��9�dy�8��A�7@�07⤀DF�Щ����ē�p��ί6����xt�(��<��@��`9��#5
,`�����$�F<�\TF���Z�k�Efd�wM})�k���g��wߣR�_�37P��)B���*$�p�K�ۻY���c���Q��?l������F��Y�[;ed}����������5�h��.����½$��?�_���^b������=�.�(/;��req��24���Q�q��t9��4��?�*��%7c�����i���<у+�i/ffn�3���i�(@w �[m���=�Ǐ���3����C����>qJ��T11�g�� ����It��U�2}T����+tc90��Ƽ:b��F�E��U/�\���x�����`��f�4�Eɓh9������˜�!������ڠI%G�PӘ����`*y� �iĥ<FdMỈJAݓ�1%�֖�Hq��M"��H����!�M����	����U��W������!Cb�T.����Q
L%s�0�߽��L�:��|C1H`:HF*�Y�bl�Q)��K�Y=�ݍ��܍?|�;pӍ�Ć\��W���?��;k�F�d����1�������㷤yy�
�V�`jzVz�x����IO�i���M��J�E� \Yd9����������J�>��-\yY?���k^�9̘��k6��ן��s+�p��[���t�c(֖��K�؟�U���D�K5���H^����/��RUQy���ʖjb4@��c�8�C����[���������l3M�t�KQ�'W�ޘG�����?����0�t����_��eA�����u��РH^W�Y��h©����X��H��Ĳ79F%7@����+���k���a�#oBg]r��u|�����z�;u�QE��(�DS&�o�d��߀�Ti��)ِ�bN���J�[\�$��˽���>c �c�$p:+$ǁ��{�.��\�pr�+5h�C�d
L��*+�T�����͒xI�L©R�1��H�i�M�L(QkAGם~&2���h�_������%�	�ͨoB���(��U�Q���)�P2?UGuy��iDc5����ǱH�It�-�c$�6��
������2�+V)�H4��T1�x    IDATj0�d�M]<I`,+��Ս�m
{Z*��"�d��2`������ouMhE�۵�TQA�$3ᙥ� ���gLC}`�2}��Ϝ�m��H{n�٥2��^�ib�E���}9��%[[���C5e��E�8#{��X�Iz�$<ũ��XzjE��{+����f֋��ҤJZT2&b��.M�����I���~��s��!-Hy�6��aF�� �B*Ʒ
N�Ɔh�6�~�����T����8�kX,�[F�d
��BWF6mR��\���L挖u�a�� �ki�@c���"�\We���顠���j9���"�>U��a19���������sӘ����h�kiA�{�� v�Z���<fg�Q�����c=P&��`�z��D=�'�P=�3�����D�#�%�A��a:	Ȭg����1�c4i"g``YBj��sCt{���9z�)�y�X��)�( $#t�	����PF؍s�q:%yMi&�ϱ�E�SR5s�b��ne+�G�ٳs�U :�܊�v��u»A����X��>e�ykT͒e�SU���^CN]gU��1�ۣv�N�Ŭ�C�r�;�r�qg4����3��R���~�{�����ċis��}�Y�����=c�d�[��o���X�V�vj��9�V/8�9�I3>�{Ӥ�9~2h����s�f
x��?�������0�x�<E���wL��}
E �|�Q�o����/��S��؎��c��5>��L2���������r�̲�lĊW�(�cq�U�*���RѤ�}8�6Vo��֓�T&���OՑ'cJ�˜I֘�*��J~��ZEf�ƭ���I"e\I��Ԩȅ,0���]1��+/���99��iC`:T���z*�b�gˠSǄT��Jy/��b���ߊ�.��9��L{���ݟ�����cc4�~�� ��6'1�S�q�е�0�I`B.�HPBE�� DrC3�`2 �z܉#_n��jӥ�Ϟ0`���/0}�-G�B�U��L��H`�8�..��k�������hu�� �G�
2k�9�s�$z���L���(�y����d E�%��
%$�.4`v1U���kw�?�2����S^;�������}�� �{���/�����_�6j���gL;�U�&�{jNXt��D��2�@� �J�F9��N��9R9�!`JIl�1�b[8|�2���k�2�#'�H)H�m���<pz����~������G���}�PFWY���˭�g�g	������ys5+.L6�q,�E{%xYd�hC=@a�C-?�����uG��Vb��Z����dFS�TB4��v������cGw��b��rg9�8�ʶ���'��LS��}��3F�$�eʲ�DJm�Ai�,g
��o�_+�z�e��@d^������TRcيP��� ��z����2�X�GL9���i�W)6��3$,4p�H�3�ѹ@)ﺌڙ�tI~VD�d&1SFV9�g0T`�ݑ`+U��:ʋs(�q��P���ҫ��k'Wv��G�v[XNS�%V��a2)/g�)0-�ð�i(C��N�9J[�4�c.6QJƲ�����&Z��DݱCz%N��Cuن�{o�`G��~%O$��` ��)��&.:S&k��U�k���{��_�wCM�2)���W��i���*a<cN�5_�Xf��œT��L~ng:��o?��kvfe�&�)PΦ������ܒ�8�ˏ[v��O`��-�*y(&:p����f���3�ރ��:44E����sg���`l�I^�}Rm�?g��y<��h����_s>qL�7ĳ���IetXXS��SY��7"z�Vc'�Ҋ�? k�_C�J�B^憛ėj!���ɳ%�h�)Ţ�"�J�3I�EQܳ�����󳘛�F�Z���L7dˮ�E,/.`~fZ�g�YLM�V��`fI�A���$�f�����-'}��i��e�7�W�?����d��g�����o�����l�:����z��:��B!� [Lt;}l��8{~������\Qc���Q�a��Q��F����L)8�RaD��J�O���^�5Ha�;{{׌ݵ֣���x!/���(Q�J�N�57�1Az�3gu��Vx�
IvõpĂf?z��ە�:����\R�L��9I,����yl�2���x%�`��m��\��E'_�z%��8��U6Ù��+���-��A�T�s�)휔68�K��ryf^��=aO�W܅�>�Y��W�{}��Es����_�V;�Mϋ���]WV/��cO�؉�8��\����3�����!'Q0BPuE�EbU�K�n^�(�)��L�]�˘�^�#`�U��=�Tw��$��9����\ƴ8;-&��R��TP�sc����f��.:�[�QMF�80���W��/�L&c˩"�dL[��@g������Au��?kJy��ۆ9���2V�x��4n#?X��w��o�u�k2^ӑJ&����i�;?�|��`����
3�@�QM��<��섈I��%/��b�$6�:�;�:c-V�+���(ƨ`�΅s8�Q[k���}x�ގ�?�ڜIl<�d� zU���[G�GO����3|�+�AWP�Lcv~�j�UER���=*zf��WE�\E�\V[t�!�A)���h�LglČ���b�g_�/|εؿwAQ�V`����X��#�6c|���ѓMD��l�>�2eS�.K�hE*{���z���58:��(��aM�����I'LGqI��F��G�8�wϹ�LU(�e!��e�n�Ffϩ�Vd��[o���`�;İX�>:܊��S1pJƔ=�:���\J��3)�=�H`P��� B.�,܎���}\whWZ�L����H1�2�tH4��6�$���VO���֎����Q.��� ������9�UK����Am��y�{	MB�F3 u��zXQxBz�����Br.O�/�iq)^0�� ���&��48�>q97�W?H!ٴ^e�B�I���jsHJQ#Hv rZT�I��$�^=�����ߵ��e���a��%V��3��
YOV��5j(-̢2?�AN���vuՖB��4?�腭6��m	���1f�Ș��=?;T+r�� ��\{��U����r]ҵ��ǸI/M�(ea�Yjas�\l�V�<ֳzx�z5>eC�0w�3�<eߥ=[�0�iH*��_����޷�J�R��?��0����Xw�M3g��D:�o��2_]{���o������G�v����!�6�D ��J���]g�%.
 wI�}��{�?7?��+3�EA���K�m=�R�"U�d�g�x�?��A2�	�+}��a����+N��� ų�&�.X|Iu�p�Xo�p�X�
x�A?�����-�$00��;�����1�����8�"�����d��ކ�ؙ3�R`���3��P���d՛De�m����H�̐*(;%'�B�X�E����%��$ �,��Cɺ�I�	8���e��JeY��ݍ��)�kT�%��,ԚC��;�<�
�5�%�Va I�1�Κ��P��A�n��n�v7¹��s�C6�fC�-�{E�<�u����L��(�,W�h"���j�fET�$W��
�dַ\g%�15
�}�*i��eg�=W=�<Fn����F�ލ��̙ܯ�B�X� 3�}��ΰf�X
eԷn n�4ْ!�]�*Z�u��H,j:�8%���ϔTfa.���x�O��g	m�+��Imt���{��/)r[�p��) Mo7޳�
�)peQH'-��U�S1�7k���.�IW�_�+^�\�����e{�uTE��=�G�����?[��|����&"??z�?v
'N����يяs����9�#�(Ago�h��sD�Dˎ1�!�dN�̕�ߔ�2~o^s���������8�}�jc@��-H,��h>3�\�S�R	�#mXC���WʨQ��ꢷ�B��K�J`�Rކ���ƉF��/	qCƴ7@�Iƴ#��8UCyvJ&�D���5��Ι2I� L�%#�{���&uI����"~�����w������}��0M찟�H�6.,�.��j�Aﳰ�ZeJ�������z��Gr�.v/U1]�c��,�"��~<p��v�q��{�?���e/�En~��
�MZ�y:`ʍ�������L���1��`n~A�x�XmTs��*�T䈐�Q�]����/G��i������I��ja�R��Y{�;_DiD��� jcz���:��ۏ��8�m�p��6��)Tg�1���r��6Z}���4���x�'�^3s�����t�t�k���?Kj6���I���A�AQ�"�� ��v�
0�5H�bK��^Jޫ\X�tc���m<���fHJuD�"��U��&��2�|(�dU�q�
�9���6���$��%� n$^g�b�F���.^�����[������i�w�j�v��v'�^�C��a���{#��C@�a�j_�6��elL��j�.;1,��]��i�1�!sk.���ai���Zeo2�\ںD�N G�~�y2"��QOn��-%�>���Q���H��װ
/⴯���3�@ma�r������~�,�Obl�?�態��,�ڍ�2S�h��T}����	�KkL������nl0�!_�����އ�&�RqW� l-��Fc��a�����T�#,��+/M�"����<�2�Awn)�X�Ғ,��)1��c�n��(���`����)Ѱ�fZ
p�
 L�L6qR@c����[)���nNT�3��ғ,W�'_eo�Mv��5Sy�dҁQ
ttLL���؈e�2�G����p,�T�ױ�O��;k�u.NY�4���+ Q7ܝ�?�{�d�%���Y���G���J}����ݩ�o38���>���|�����y��V��j�y7�1ƞ��r��D�¾�_S� ����n�-a!�kB���ۈ;�W��m�&��̞Ÿ�$PF�p	@,;f����<i򯹇T�%���3u3*]����1{)��3T��h"g�,g|����Hg�&1gnǒ����|<	�-h�*���.�P͑l��+���9�Dl/M���dƩ�$aX�y�!�� Q�Hl%(��OδqQ�Ҍ=��G� �*��ZQu����u�&�Nmеo��r~j��3���|I��pf��uʼ���^5+�5�� 4,���gtq�8+�ć�^���<��YAR 1f�8�~=����i�E�r�5a3���-5��xlmM���ԟ��֠��"��$��¯ӷbhðqC"m�}Cm�={��*T��9��֮4�����	��"�ږW
�ͷE���$n{0ϼ��#��.�~�-d�l��+��-ϺϺ�j�^����,f���$��|Su: �����bc��G�8������s�h�D		��+��n��Q��3W	t��z��	������Y&Cj�2����X 7Y��y��s�t㸗��C2H��hP�		��R)/S~݁)c�f+eT	��=�϶'��Ѐ)՗" �u�끧+	 ʉ��#aL{L��^"Jf�x��R����G4�S`J��a�b�Ea��s��~���>LC���92�[#�/���6GuDd�D~c,�UY%�1Au�H�9��YXS[�"�0�Z��SU��튵�����po�����\�����p�u�x�އSǟ��?~�W��W�h��f�����pa���Kn~t�T��Ώ�_Ѡ�B�2�"/���^�������l���=r��o��f����h����e�� ��赛��ۤ�Q)�P/�8[���
��?���U��T�x0-/,�F7�R����I.�/|����W�{�=�F�+���`�^��ku+U�h�,�\k��J>�D�X�cx�.�:�f$2�nkQ��/-��b�|�=x�|/�8�O6���"b���qZ��4�vz};����\Ó綱5(����.`EMx�ښ��

�Je~^���^�d�V閙�c0�m'Sa��\�>JI������y�17S����c��V7����x��p�B�Q	O�k��g�ƞ�HF��}E��q��M��'J5c �?��cm���-�!��4ρ�/[K�gxN��C"�3��+���lO��6JT��-�g+�>$�����ك%�d�9��y����~
�A�8P0'Ur1@ʡ0b��9l^��B����{Q[^V`JbՊjU'��QB�BQ� ��MC�g�Ֆ絒W̡O�\DB��ǘ�I�6Ĩ��|̢����ݓ�2�ٕ
�S2ϔ�\��B��4����d(���n�a��B4����A�3Ig=e�3��(�,���F�l_�+~��B����w��̛�~���Z�g���+4��韥g�M�l����yyb$��%��r�'�Vp1�i����g6ɨd�y�����LM�?Ld�hA,���+�k�4�xV��w��C��z��Dyna��+k<1	��)����*V�)��$K�7.6�AM�]
�lt6֤���4�doe��@��b|�v����gصj����������V+`(�v:^��g��#��^h(�9�Q�`ٖHW�J��<woηh*mԱ+�/Qgd?�$�kC�mE�ee!�瀗�:}����衩�:��X$J:�.�ɋx6��?�e���,����ƫjD�M���m�p���/�����y�!�32��"������r<z���<$t����ʀ���T~%Mw����I��9}V�D���%���)�R+$xQN�m����c'8�O��xiߧ�͙Q[g֦ ߒz��O8T�8f��g�T�0��٨�{"�YX��U�H��̇V���_�~]�{�8a{�8�炔5�5Z�V��-T:���C눻��W�wLhy�I�~R۟i��~��(�c%�R]��-���y�p�Pj���Q���X�٩2f�����e�l�.�Z������(@������������F�~�eFd0yV�t(a�d� )�bE���H@J��ڟ�p�e���X�R�9�i5h}ς��Ȫ�����H�|c�(B��Iqi��|��Ts�k�Q�%#g$ò�&CT9̔��Q!��cJ�)�d�jU��4-���C�I���2B	���&�vO�0��
*3�����Yb�S\�|^����6��r�c�9���x�n��ӝ��������w~T��Ƹ�A��D2<�,��YaL��q��ά��:��u�6P=��)�&���6jt�l]�l��?�������z�����3��'ԫ%����xݫ_,��_7=�f~I�S\��o����_} ���Je�FM�t��{���g��b��k��Q@G����gp�#Љ�Д���	ވ��×�a~��� B{{�6���8�g��U,��13SE�^A�Z��Դ�jr�)Y��kh����	�eeu5��|oM�U�����$
Q��h��l�d�F���l�_��sFD@�DA0N�A�QQ�QFA�n��;O߳����S�|��O�Muս����k��n��c���I��~��o]r%����cv�����G���r�]Z������E�<�B������96�1u�|w�k-a�t[�˘�ce~?��<�'�5�r�زI�i K9�8,���-wp�U7�����[EkP�L��l�[�U�?W3�h�PA�_B�6���`��%�8��n��
F+��V�P��719���� Nz��d�9����˂_cat~�����q�}���憻p��/��ґX	B������(�LHVm�O.1s��%:6[6�NU^����O�k�#�}���̪�>��]����������M�k�g_�ٽ�O��.M�Ҟ� �x��cJi	+�u���j�|�.�(��b���}�0�w�f�N����(g�e :�k�L+�>�sKh�/Xe�IH����(�W�C��FeVd�l��${L�6�h�-"����ag���~R���c��*b%U�$Z}�^]Q��	��^��]��9��n��M�Y��2\���˷�ۦ:��!�`����ɬ������֛%O��(QȎ���    IDATp ���w7�\�rH8���l���I��Joڑd��6K�l|���?���2q���Bb�z���뵉Y�^9��3�9i�:��甪�*���D���q��8��xQ�~(�ZJ$$f-Z\���h:���լm�밅 �A�� 5֤�ΐ�\� �ɺ�8���<$�Ⱥ9M��z�ȱ����S�>S�j�(;��Ԁ�U�D���Q��'��4c��T��W�x]$0S!�S�;�ȹ���jGHq�U���Ň��OG%�%��1�cU����i\T�"x�51��b�p�T�եn�QY�gv�29lC$�	R��������Y�����_�:�֫��j([���2+�i���/��
`����:y��A�npd�sD/��9cJ�dAh�L3=�F�jtӝ�`�9�Nl�3'�I8ϑ�9|�GE46c
��^~{W�]��G�(�ϛ�#}i҃�qЌ-���?Vr���$��'32d�Yܒ�k}��w{��'\��l�h@�lR��q8���o��+�3̥�rbL�Q�ch�Uݕ���~v�?% ���0��xÌY�-;�	^A%�C"�=��Q��LGY\�p1���+��꼵Q����.��k�Pi ��T���UJ��l�f��M]�k~4���+ѐ����9��l&_>]�#�(#kw'[�d�j6Z4���E�$U��&+�$�+%���GG0�{���:�-=T�cZB�{r����
z���~�h���hD�S��sr�����vV\[m,/,�Uo0��� P*������uXH[�̕�r9%|�|.��9�X��2G;��IbRLO��'��g�b��b
#J 5�Ql�%O���t!��ÚK��(I"�G��:���@h��E�}�p�a�d��j��w~�3?��2��O��K^�G�`�҉̡�G��8����~���A�?��ft�E�ANNM��ZĦ�
������O܊�T=��y�7|�_/�/n؋�F�Z�^[� ����]���x���?"�^XY��w�[o�#�މǜ�pL�gc�TF��$�+tu`��7��^�������U�mo�;<�GIW�ybl�>�7�[���"r�*ʍ��D�d�K�a��)��� 1@ο~5���I���:p��Wcl��'<�1�qߦgW��3�.t^�����{�w�k_˭��W������?8	;b����p퍿��ޅް��S�֥�Z/��IV�ˠ�nk[gF񼧝��ގ��2�+˸�[�<��|��q��i���87G⟭���V�����^w7��՝����Z'�����(�����G���:���nܹk+-��̪3g�E�E0�TiD �0����M�
ZA�]q�"�?oN��0�;��`�)i]�X��;��:j�bLZG2��©$[&���Q��QQ�I�H�� MK}���� �@)I�~OS����5Ln:L�������]����.���
��dG6N۸�\��tJZ?0�o5���Fҙ���@��.l>?�
��TP�a��1a�D3 �5�.����d��ɍ.z�&��ʴ~�ꏁٴg�kF��iy�$V��3�����J$]�f9�orOT4jI
��x[\�$�Gɣ4z�#�8	H��G3?�pdl��k$�~_t�
��H��1Ȗ�&�Ai����@8b��(9�$Q	��$sQ�uQY�*v�p����I��8�����9��k8��l��1g
�:I�w�yRj#%3�s�Bʧ}�D@�*[�θv�IT"�K�~:F�[�pV��b�5AXBf���'@Ir�dzI����cơC�g��⥫�{R�8��Q�=k>#K��o.?ڢ�U����F�xo_&��8�$�0"�h�g�IߔC�"���[���H���<�	�8�T��&��/(b�ˉ���3[+T:�WQ�-uy�^IO�Ǌ�A3<�g��v���ǲ賲J%��J�tT�}"��f+A��������؃�J�K]fn�p1Z*(ݭ�W��}7+F�D ��AL�y��|��rP{z^	ScD��խ�C� ٗZR����c�x?�����,��d�U���(! 3)Z�����7�b��-�{N����c !6��H�k{�\�	�m�(d]&�r[k-*��%P2����* ~�h��&��v��0I�.����B��s:�T`1bG�ؚ��"��/�^1��J����*����H�H4"O��=�|��)g�,*ѡmkC����?%{%i��*�%���&�&�b��e�Ӗ�&P�?>��)]~�>L�x���aUJy�%T�Cs���j]��}��=ő���Z�f{��2���b�8��\KѼZB� ��W�E����x�_.5*��"B�-S�bw;�p�_�w����FŔ�����fR^VL�0����X�`ۗ,�7�zL#�P:g��i�-J2����w�+ȵW�o-�M|��w����c�s���?�g�<G��-o�[��K�����u���t��p�.�ҙm����|�3��?��^SS�Ѩ��������O|�&�s6��<�>t�Wq�틨�J��֔��]�-�U��?�x��o��m�1�qm�l���z<�aG���7�B+�`��,奺�2,$x���;���6.���Ҋo�,��{�k���?\�L�m ����8��oa�YD�<�Z�fHF(Xt���I���Wʵ�qb������G���վo�����aG�2}b�}G)|�g�#k�	|���q�7~�����jG����g��w��=a#FJ�|�:�O�ه�Ͽ{Ҥ��V�ڈ��pn�.+��l4P�7�?���'����Ņ���q�/�Ƌ^�l��9y��`K�K_*.��J���]��U7�����f���Z	/}�3�?�#lٜCg �] .��z|�{W�7g�����f�9f��a΃ �"�o?	-0��'K��@k�H�ޘ(%�Hj���ٚ
E��YrR�(�~�=Ӊ����+�0�,��0Aer��3ٿ�\$�i��1]ٷO��R��-(OM	�rn�U$��U�i5�>��hAR^KJ�Gk�N��W��y��"�r	1_O�j��-�њ_Ԭ0��K4�[�[2�%UbA9/�����b�8I��VqR�g��� �f����{������B�gP%�P����Ҥ,_c7�{�����MV��yb�Tug��q��4C������T��>��F�,�L��� Y)��>��cZ��5���*�9��;0JR;w�t��ɨ�C�Gd����k
����*6Yu}*�"e��I�B%&�ߣ��
�M�rwp�����Y'ݲ�L��#��&L��5�������J*��3� eM��8�/\U�(��6�׉5'gRy��U��������	���X*O��d���1�E���0�ʌ�XL�\p���<��ɻ��I*9���p�d���U;u�%a���T� ��ٗ�����|=��T��G�e������;r�v&�դD�1���7�#��\�%�G _��8��
��/�F�����&*����6;&C&��l�%KFI���֢'�.���ۄ�<��z>#�3����@�q_��sP��3�Nv0MbR"��V���ge���_� 
hf�<́:�U.%�!ʌ�ܡ�����A��z�S��٘lUy�Q��*�H
	y�S�X��=�'gj�C|�&f|��R��[�2.��]N��':T�ב���ތџ�I����B�����dڹ�� n�F'��z�LڪD�g�� ��\��,�(�Q�����b5������L�4��!0��YbuԤ�t�՟��6C>>'�)�N��T��>��wݡ�iR�k4��=����]��}^)�4>����t����C�vL'J%�9�w���������(���LE�fi�$5�W\s4��� �����S���
����T��nޮ%R�g�I�0����_~;+�������q��^�㷏b�����bZ�4?�+�e��s�:���2���LE���LE�y����G*���_M^g������"��y;�8b���p
v�d*�m��ߺ�>�lIk������"�(���L��F�Ãs}|�������ڭ<z�!�M�aei?�9r
��[���ڂr��)Y[$0�a����a�YD�Bg^:�RB��Xy��?����W>[',�2w�[���	N<�Xs�N�眠�TtF��ʽ��?�j�-�}}\�?��.�1��mo�+���=�2�=sh8����/~��"F'6b��);`�,��8��,���65�g?�w��t
8p`����裏��(�ײ|^�Ua�+��e?�_��{������ᯏ'<����߄�S$��C৿z����x�@�~�긜�y��R��QG��Bn���x����W�;�Kv������񰣎��[U��L��E���G�!pp��5���+~�;�ލťU�:ml�2�w��5x�����2���'{�3��fo�!����^#�K�=x+�n�t*3���}�$S�b���
�G��=X��3�� S���2C K�Y-U�&h�\^wtc$�[�I�N0� Kn�##�NM
���XqI&i����0��bu�~,8���7� Ӑ��z���(BҔ�����g�e~D�������c:L�{�ƚd\��zЭ���͎�$�e��&�
�5)�)q�)���`3r֪-Jv\+@�~Sbd���K����o����*Ӷ��.+��Eb��k���\�%s��f�f$2Cp��?�Bᇻ%
�{m/ZJ�Y�!�2  ��ſ�IV������\��H�E@��"'�D(�6^��X�!ՋD�+�$V�+������y���`����.�
 RQm� @n�T�b�JM��0M+I��H��G�C��Z3� �&�O��@�3�lk`1*���N�O���31t���%��?Տ����[N�� ֗j��w��83?n|�XB�҄;���-ԿE��k��������DD&)V�3Zc�'fl.�uE�}_J�=�������5!�$[V�5�05�}�C��`�qf��xH2������I�p�J�L�tH8�g�6!~���Gc~���z�u=�,`�Ҍ@��Q�Q:�����������<��"鑵��̿\L-֤q)ݴk���a�05]N�%��6u"[�u?��.�hHI� �2xϞ��''3P}wp]��D�S�)\��%=���:��StB����?��:1�u��m�&}�q^�K d�N����o�'�7�9�-�;d�N�*���k���{dc�!�h<��ag_�����UGճh ��.���JL��ڐ��<I/u�W>�c�xVZ~����F�H%e��%:���"�)��"�$����1���ֈ����.�$@K��>D�1�7@��Q���n� a6�Q��/K�+yj��������m�=���X����զ~�����ȕ�26.w]Sɐ3؀ϖ3�+�&�%0���WӲzLL��Ɉ{��
a�k�)��3㟼�]�{u���11��v��F�,M!~�o9S3?�
�_{�zU�
US5ć���)�w�T�8����]�b37 q�����ige���7gqԦ*.���b��ZRi䜭o~��8����Û��7x�_�	Fi=�ɕ�iB��S��U���b�i�3Ϲ_�֏�j1����V}��������lGI��y���]��O��5\�,�]D@iNy��̵���>��w�������o�s���xؑG���G>�(L�73&Ҳ�6��Nw���U�.4p`������w�_�?��Wh�pĎ	���^��x�Q)rb^���_����7���Ǻ�-����^�d�y�޻�ZG��Ű���7���O��NW0�a����ko�#�Hu��0G�K0tV}%���?��=�;x�EI��>�����#|=���v8�2��O�} ��2�v�*z�
F�֣V�:3E;oL��鸣YrKؼ>�������u�#�$X\l�?��\�����b���$��e"X��A8Hyv��_\'�����{�g�,��:��ر	�~����?8J�x/	L��i���9Xj�����)Uj��id�� ��0���o.�W{%����p�װl�	n`��tp����еf�LF?�ɐ��@��P�'�U�_�{_�Yn;��:X-��U�Dk5�X1%�esL�脓�*�6sڤ�{�`��\LK��2?
`��\TC`Z�М�Gs~�n�rYR^�-���Nu$48�;�ɻn#k8O�r�����..�Y4A���%��ba�Y�H֛�V5JfH�T�U�ڵ�稚�aD��"U#�r�d�4B�	�1�^�r���*Gm���5����=щDa�e��-�2�V�˝dSЙ:�Zb�&M�hD��g��t��D%�F� $��y_;ɼH4�O�.���d@o�|�}�z/U��$��ꚳ���D��^I��i�^�Q��K�C��B�����*s�g�EL`���"�<9������AB��U>�cQѴ��ϻ��Z�l�7�b��Nr�{z^�f&��~_�aX��9\�x����0f~N-z�i:AȺB{E��û�ʥ��7�k��ɥ�3"#���JX��-=���t����� ��H�[Teq�}_sI� �Ϩ8��ΐ�;q(#b-;�6O 4���G���`NfEv�/��ZC^�L��R�N�{#����Jr�0�͐�J���I�df=�[���٘Y���g��
�5��' !>�萴���9��%��NFioeZ�$��^���KM�Rá�R����ED�����)���3WM�����쁤��+���-v;�t3���G[��'�����tiz���S�s�2 ����q�?�ΥhI*�ih4y��ݑ��Z�Y���]$�ǧ�ب�_�ڟ��dZN�,�3�y�)���G\��<��g`;�d��=Y�'��s7��ʋ���g��Jʙ��GJ��)�}D�&F�?�<&(�%�hJ A)��h�� �l�X$%�W��I�3�a�,A)ի$FL���bZ��z8J#�1m�e\�kw�i�,�`�bF�ȱ�F��rK[lQ`ZB`�W&���h�4��*���P�#S�S^1�Ok�1u��aʷX=�����M��0��p鿃p\e��=��_�?��U�Χ�49,9"�ADM�^�Q��[u+9g\J��8���Ķ��.�i� ��2��|���8bƥ�_�c�q�yb
�����X�\����@��,0��G����\��W��ϟ�t�et;T�E��8���ގ'>f�w�	9���9������i��ҩs��p��u����<�����u^�p�o����.�ԺIL��`�֍ظa�rQø�Fkh6r��_\ť߽R�}��\�ޭ�������2��mŻ��j���'�\�]s+��Kn�i_�:fX7y&&�U!6Y��UK�$�
$��|wGo��O������������/ú���<��2�D��Q�Xi��hw�on	7�zn��A\�_�a��E���Q-���g?��1^�Hb{���?�g��}��`����'Qa�� �%}L��mn�Ě��7�%^��c��{�Ud�+m\~����;��g<�<�x=S�����;6�m����&�}�!�v�صw	�Zxh��f�v�-�Kؾu���ĳ�|�����B?�� ���Rs=��\C� F}GLvؘ�4!NC��',�*I��YrɎ*��"��D)e�jv�s��`%� /I�U;���!~0��Hi�q����]wi��K��1�aC�\+Y�x����� �'e����CX��G�:��)�i[3C��5Z��J`3��3Q�И�CwiE�\�ɬ����.�����&E	s���졪7�Y\F��E�R)��(��a�7fG	y�tP���*�}�^��%$jnn`2����{t��A�ήzA��(;1�x5R�[}��������%: ��,��T���T�.��̈���Y�M��l���'迻/SM��up�U��P�V�\�O�Y����[�I�uzLR$�yT��J՜��e�]{��ⲽ�)]��֐��d���'�.@d��%�Β�@w�.ӎb{}U��5�ȧ�@��I%՝<.��g��+=�׮    IDAT�9fv���̴=a���'��-�$�	���*ک�OW���L��0B��	��eX� u��������۠����H���Fq*e�n��n�U�,����=K�6���~Z�����;H^?=�ٻ�2>���ݔ5t�k%��J{��g����{�$�1J�(YG�Q�N���P�\N�iV�Z�����@�Ÿo~��Ʀ0q�ʴ�1-�O��L������₟�!�O�0�2������I��l���N�Cj?ar� 
ܓ�[�2*TN�d���-"�D��!�z�g؃kB�L�� q|3��I�$�&�6FL(������2���&�Y��d?[���]3�)�1g4�R{�I� `�=�A�g��Lf��5��^#V�J������N���<'K���� �+��Rr��;^�H��������\�I;�9�2�D����r]Jxs�q�9͈)�N��B�&H���=��2*P�����Ҝ��F�M_�m�"O#%Ʌ	zke��%�!}��Q�Q��E�7+�jn(W^��k7Z�6ţ/`ZQ�t�16�I�������*���./-�۶�)%Ĕ��I���-)��;�t
� 6�Ry0c$�jw��v�N;�u8q�zL�	��_�U�.p�?�����*:Ś�u��%�n+�X���2~]CI���Z�0���z+�(���#�p������'�f�sɥW��}E,ԫ��Ex���clRt١�pGp����PL�]��\�O~�\��v0Q�P���ۆ�~���= ��ýs�Gϸ��� �(��v�{�+u�/x������	ʕmK�}�C8��/`��i��m�Z��3�2Ob_��329�@�������Xm�Q[�A�����'������6�es�z��g��J�u��<.��F������b�L�4��\��LL�KV��ݨc�Y�öW�o�y���|�?���}�h��xғ���۷bf�]sH[����o�A�����8�����.n��>��^Yt�Ky��3���>�vL�Pr��%/0�ßߍ3���{�i��)��z�d�uw�M�Z����U1��g�q���$Ǿ�k_�w/��w,N:��P��1{`��s��.|e��B�"��~���"V������އVsU}�������h�r͋j�
��m���w����8:�*J�QT�#ȗ�C=�IRi�A�4㏺���K��H.��7�#N�d���#cA�n��V��0ٳyvV�qI��Ě�ʤ���>���!�ɢ�L��1�@��M����iIz��:v�6k�8ȡ�qG��`��27�jm<��G�'��1x�Z����-ݗ��\y�4x���d��4��zMpyht�hM��)�Or���f[sMs�6
��^�s(Y�)�-#�*>��
b1�nf����=�z��);�tГ�uɋy0+3ظ���d>n&`ɲ݋�oF��H��ۂu��Ck����W�yv)I�ya����JY>�6I	�4ڒ	@㽗��1k�7o'p�j�P����J�}�����
bw#�[	4o��'��C�[IO����2�>��M���0�ɨ��G�O��Y��5D�%��L �U�-����IzL3���]bg2�I|E�٠!��!U�}�ٽ�^�0����D��Λk2?���)X���]����������&�F���@&�YBְ�׊�I���p��Z� Ie��q��6zĤ�!L��i��?$�6��~a�3f/�B ������k?o}��\e�XHH
�<e	�4����>��*�ޠ⽧��$L㠈�80������f=AV��E7��9�Y0�}���d�An�SV�4!Fla�_M�_�~̂>h�$Fx��>�01��5�q�a�$�Q����`�Ӯ-UUٿ�~�����g\Rj�Ϯ��F�%Ƽx�N������F�ٽp�7���,�j��4W���E��s2#�:�B���YKr�~/Y�qgL9�R���֏8S����zO���x]}t?�c/F�'�&�Y�a�d�Fg��e�&�OR*'J��:/ē�ϒ(����?���[��էS�d4�"{H�}��'�s�{lT[A2��P����Z�`:��a`t�����*g�̣�`�W�"m�`��A�����~1�c���(�]��n�'p���u�yK(�Ԑ�q��q�j�����O��ǔSf��Z�1������:��|�i2�i#�2��?�Ϝ�:�����&h�t]�>\��m��������.瘆�(hd��J\B��?��ݝ7�ѣ_F<�k$ֽ���`u��A���p�����U"�0���ҫ��G���+�������L���2:֜fs2Q�KOrx�43��șbJJenb��tb��7�<��Ljh���k��Gl�G>�v<���P��D��L/µ�����rԜ[�4��&F�-���� o���0�\����}G~$6NOcfj
�S�2$�Ti�����OG���U�i�U�m�k߼߹�*,./b�acx�[�/x�cP*v�G�a|�*��{X?�㪘ZU�͇�&h�h79�x�����ߏ#f�b�_{����K.P�a��}r f�b�
+>P+++j�����X7�	��:�p�]���.��s��g>����'�c�Lʛ���⧿Q��-��N��\6gU��P*��m6V$=�8�ǻ��2���aL�7-��u��^xڻ;��s�6�=��������$�'֡\�btlB=�#c�P�T�B���G?�%�� �v����(>p���g��R�2����w4��w~��8:A�P���\��亷��Z�&v�:{�4I�쨌
�����̀�9���(y��д�\&b}A�%V-��1��$_Ρ������HV�\l��ݶ�*
�05��$Č���I��uU94P�Cƌ ��Y^?���0�T���[��F�߫p˯x�U�b��`��p��`���,z��(�����;>�����xIg'����U�N֙sF93,��`�\Ǡ�B^ �F�hx�z)
��W�:�rղ��YU������y�����X%a߈�
K.8���1��{T�T��9��oJ���蛼��|��:VZ���GEȸ'�f=v��
�o	���9�h��I�'S	5y�]��jٵ���+VIR��W�����ˋDP��v_�Q5�'��������g��������W��O�+#�U�d�� z
�dy���q�n��5f>����I�և'�z�qVe�I�L�٬�!��&Y�_�Tb�o!� c��>gHu�bs"�3��`{����|+���w��D"�&1n�C�4�%�v_3�Q̗���r��X�A@δjRZ!5�r>cY��A��9�h���l����Ur�O�=� *���,������(�u��P[�k6�L�l������j|鸉Y��d��L?b����"0�\�@Z8�Q_��ȁLE��wHy�	;H���ڂ�ua9�UN��ȏĘ'U[X�|�ǌC�{dƗ1�M��6�'��#C�aO��QN��}��	�&�LF]�GI��;�b��D�l����F�1��Z����M
��9�Z;R`��T���d�4	R�+�F �g4j�+�����[�����&*�Y�l����������Ρ���P{�Z�'�{��IU�g�Jn��x�aG�1%��T��y�K�%�~?�^��;@���W�̎5�����!$Y��(;V.	L��RJ)/�)�E�U��+��jL�S��I��5���]�d���>��Y\�{�͊cgF�< ̄����F{H�H�W-�+�d�D��i��i��������wFa����VN�g ����jO��l�bڡĘ��R����}����ᙩ[����X�d��@�����q��ހGn��P������px�	|�+W�[���̏�3�Q�O�łX p*��?c�����ͣ�| ���8��q�g߇-S�##'Wދ/�	>{����������U�Rlݼ޻�f�����R`9��#Q`�J�Q�������if6��rE�%�x�o����ŗ�z)���N���7[趗q±[���;��Զ{8�N��7qӝsXnPfōs�8�r�ĺR/����k_�G��J������`ff�##ƀ3V!�F�גV�*��N������q~{�ع}�x����b�t ���0��^|>y�E�[b��6�����]z%7e��Z�e�{�8��1����a��I&Y^i��[���¢*.ss�ػo�WV|�YA�h�ժ>׶m[p��M�k��Tq�o���SN�O~�6ۓ��h���az��<+D��*��]y;�:�r��G���&�P.���pe�v��Vc��<6�vq�_�?�8�1N89Ro�p饗��z�cO�����;�6���Ԫ%��Ɇy��jh��u��g��2n��LM���~3^��'�R0�{�L��1����
�VP��}Q��>2Q:�2�x��&��^�е �BKR�Z)�ę�����5C
�����~�%�'[ffp)�0 ��8�YU��Ò��`�'���9^~�ZAer�flIڛ���*X��K-`�ic����� )ﺙͨNo��܀\���ӹ�Ī�p���YVW����>o���#>A���U��G!�a}�zM�{|>�>��6��&���*���t�S�f�`m����C��!�Y�k��=f*^m bk,M�F�E��%+��T8#��,�G>�h����I	��5�:2V�tz�P'��?Ѥ*��em	z�0�C��f�3dH�x��V�D�ADV���վ��T�"��&���kf�`Å�%�BaF�(q�YW���0GT˨L��$C��QI$xz[�EʻCf�Ij�)Ht�Y䘿�E4x�J}W.7�~B_^%�;�����,�uS���Ҟ]�k8$N76�3u�L�J�{�PI�P\�;�r\���k���4���l�+�	V,3Se�஦�nꄂ���|YP	�u�ӴZj�X޶`?,�<�{�����+�Zw�@d2���&{�+���Z�^yZ�<z�R����R�w�Ϋ�w��\>ֲ!g�^��#Q�_Y���O������4��jT˽Bg^Nc�g2ˤ��UH�����!��dq��L���ʝ:��#,f��ˬ�g��I���0�-q/�Bf�
��)mT��I)~�����%Toϓ�*K��:�9���&�^�� K����L���ӄ�K	;_ݔ�%�~�^u"1Ƞ����I���KU�<Ǖ��>�J����X�E<��2�D�\^�O�~��}/x����B�ok99���������@<� "��b�~�|�D��������,�t�G_�5�k)Vhi$���q �<}&��R��NO
S���k<��R*��&'&�$�V.�A�������J[�n�L{�>�=>�r4G�V%A�XW�0e����#�,�L����_����X�Ҥ0��y�Tqf|+8�'B�'W^���������m� ����]>q������⠊v�bɧe�Ɗ�a�f�7�pW[��p����e�������;�,���X9 `z���骐�`�G���w.�	N���X���+_�B��o�;�M#�g�=������`���غc�1^��=���{pםw��G=�6 Wb�4'��Nx�@���^��kp���b�C��c��>H`�ÌQ0+�w�g~��~�2f�����	|wZu�+�5�'�~<^��L�fa�4�ZH��5�L��Z�dÙL����� ������G���~};�:r3���W�E�y*š\��p��K���O� �Ln؁��i�~`E���1��Kv���#���3ߋ�r�eb��� �6�mL\��Rj}�Z��E2��6�JZ&C ZX��3/��x��.��)'��/��M3U�i�+`�|��[%�}�@�|��Q*��(��'���*��%Ӎ�=���W�EO7)�����!v�ڭ��f�-�O�[�v�x�L�7�,h���{p������ހ����w��{�P�[R{���w4��w�b:a�b��q� H�3�DE/���qh�=$&�Ie:v�<d��d
�J)�~�Z��?�S;�������}mN�pd�h��l�V�O�:�q6.#�w�w�&bҜ\r��`0޼vV�ِ_�\��XMfH|��4�x�[�b��ma�S�Ll؄��a�/4d5J�(��8m/,����
���"�IVJ���I��.t��q��ɬ���ژpp�h�+p�VEV�\��J}\O��zji�DY���"��a��m�Z�a�	���r��!�<�zU�9�!ӊ���y������=���Ԓ�c�A�݇����D:�q�
GT�\B	K�� <J�,�Lb��
uL��6�V�[��U=�N�O*"	"����E�De��ٶ��*E��~K�&Gh�U�mϦ}ԑ�݁��-{C��Y��ǥ�cs��$��+Uݝ6!yu!�6]ʩ���r��&�Lk�ڂXp�f��>� ���u�XK�L�aI�	Y�� M6Ds����LM+���T����b����C~�C �2�������.k�CO�ǣ�5�T���۱3�/�
;	��U�2Yu�o��0I����+��c�~��H4�ZKE��<��-��d^1/f�:�p�O�f��q���wM��9��uFd$�����\�[��=�dݥE�X\O@~�N�H��Z)�����<O�f�E`gz�=��.�u�b����
�.Q��+j����"y�|Ό�2p��1OTB�y��߳�/ٱ�s�4$�	1��0�{�_=}�����kgx���@X1��URŶ*��UTgI�xEV@�[9�z�9�~O��n����ٲ���qY}*��6B�}�x�N�HI$������z��A2!��R<���aİ ��h�g�"Fe1k�ݐK�e����+����n!��3�2��#��E�{�q�J���)�d��I�kd��n^w�М�j����!sJ�-r�6�Ȃ� �r����g�hJ�K�#mA�,Ӥ"]}	t�ٵ���{T*�/\��`����
�-������
��P�K�o��3��
M�I�Ƭ�&���\g]��y�n�3���ŀ���k9�d����ឥ!>y��p�o�aqH�4�� �He��<���PiZ2V4�5w�q%�k�^��+o �/����2��o��8���`a~�x������8|�
9&�����lONN�L�?l-1����}_7��ȸϨ��{� . W��V\p���_߄���;q���JML�>{�e�kWKM�#+�b�m70l/c4Wǟ?��w�d���<���7�'!{J6����\��d�@a����:�^w�\r�����E�y<g��3�H�K��'��*��%ӑ�IUL%f)����:0�fq�ѓ8���j�?��R�dF��5#��H(���5׾�'P�j$�����Ň��g����S��x�s�ǰy��E�1-�����V�t��WL+#v�����<:�:�y�[s�8��{��j�Qg�L�t���([�{��!u������λ�i�����a������Oy�>߇$�/nk���������r�
F��!_p ��X"b�p���L�\v�y�~����!F*�)`�X���X7^U�V�|V(Ͷ�������hw�7��7{h��K�Y�#�f �L|,zk6�a>k�M?v�%���C
=�2jS�1��U1��x&6J��8�b��w7VU1��Auzm&�������!� �d"^�R�����%W�uɾO��)M�!?:�/V��� ��K��a5��H4��i��l#Wo"��ڀh���Ǫ��J��;�9�N�aR���@��)1��8�l3sHg�E*�9#c��o1%X���0Ǳ_=���a�LN<�����H��E�`��Y�� C�KA3�s-[��錶@���zHe���(kN�b����� �ؿ&��ٜ>* ��خ�*Ë�蓼JR�YĂ01�o�Ry3ِtZ/Q�q��Z^d`ϓkK�=q�$פ�1� ��G|�����5�ˆ��O��c�Z$�����p�"�^�Z���{4�u���k/%BҞ3���q�`��BG�_}�ILN���    IDATd��c�����L������}i<7HXY���8�j�A��'�ٳ�*�Q}L�� ���R�N�=��O��c-p
O�jZ�6�$2�������7�=���D{&��ҹȉt36FB���گɍ�bY���ϴ-X������rr(#�M�Z����Uk���sK(WcA3���=�|��]J��i��`�-r�O�Ar�T�7 ����-��eߟ+Q.ߎ��KW|'y��t��?�bQ;P�����j$f���!�ڇ�~�Q�=+�� �
��h�o�'vz�r�O	
��}��R���jj?�}�?�Ks�,F�4��Q�O�c�㔱�i_���b3�5�=!F�g+����M<e��k��(�<��=�r�W�iĻN3���2����p{c�G�UbH����ݾ )���N�J¦��3�&K�JD~��BSՔ#� �Gcd�/�t�!��*4�d��J�6�+u�[]t	GF�Q�eƎ���5-D��O�l�l�W��h��*�屑0�j�W�)�`JB!qJw��Ѐi�5�#�g����T���=�������{?�{et
�ĥ2�8�K_4b;Y�}�$���ۜz�A���A��~؋��^<�[p��ǎ�Q-�e~�_�SO=+����?{6��/��;7X�)�?;݄)�i�d���� ���ES��w�]�?��A���/���ã�݆�}�8鸝����O)�o����vO�u�̪��i�`��������>SUz�L�k�&,��|���7?c= Y����ް�~�p�-��aG��[��Z��y��>�C��K��GO�����_?cU2O^T���Q��
�+�@{'3��>�^lY��q��LG�e����̬�qv)��gN�w�v���\�cw����a�Le7�Y�ߺ�&|��b�V�7��~>�����R�U�W��0��䷾/y�	0et��`�27x2�--��ex�<"dq� �v�C�ԩ�Ǖ�y�m߈SN9O}2{L4R�{�-���?�vn�~�J��1S�*B��TjFڂ�#�J��4`�!���֊�֍`��f�Gq���ذ~������v�����!V�-�?�����.�1�T��J�^�VjGh U����#Qq #@ܿ���SK�,)��3t�q*���ȏV�;���Bf��6	�\����{P0���4j��Cs�W/�J��z�kt���@���_���<��c(�� �5�i �r��Pvj,a����d���^m�=rI��J��?o�����T�ɕ3�*�d�Y1�p$����)F=�U>�_��&^V��v	��K��D?����$�R�#�^=�|`
�z�j̙��7"��Px������<��,� z�4�9)C�+��0Ë
����y����ɽ�Xꮊ<e:2ED��yR#�����q��/w�Ld�QMwF݀i��%����COb�K�J����=����A���	� ��/�z�R"� �L�'E�$�^[щ�0�$yk֚�.�"A�\��7��h^G�� �m��R���z?n��>�ʚ�?�bm)QM*��%�^N�DT{�Y��I_{>[]L�J	�9Q�w뙋+O�}�4bJ|�-�R�s�\��R����}���)���Z|eA���ɫݖ�<ӓ���$c��j����I���5�B���^p�טE����)�w)Y���}��b�:S��0Lϼ��@$�.{�;�U��z�H�x�����R����������t�'�+Z>O6"t��l� 9�C<�z���/�"����e�k���Uq�����p�X%��I?�Z�&�RB��Q{W�_�ʝ����8Qc��Ee�?��]Cj�f�<�+H��[u#־�;W<�2�������T�w_��g�޲�w~�:Qk���7�͢i�D��^�$G�(՗��@�4՘��4��
>s�8���C���*�����X��VJ��V���AǑ0�J����bQ���&/��k=Ɋ[�͔��|�S�)n���@c��6߿REi��}�$�nT��Ӥ	V<�<���V&VL	L��j�6ʘ�6�ۥ��R`���
�7�F��鮢ԞǑ�s8�o�#6W�J����p8��`���wqݽ�XF�B�g�����8���8���c�~�����4�S�U*����<���W��1�l�yg���F@�!ӟF��+q�i�aei/y�S��7�;Y1�ï/�C(&=��i摟rL�Cs�Y~���p���m�܄G�y�����7i��; 9�"ܽ���F^cM(���Z@gc�:^��'�5��X_�ϫ�9>�R�~�E1 �[�'��m2
��&�B�˯�O�q��2�9�-x������/��jy\����O����"&�w���%�D[ <9�;m�k6V�kģ��Ɨ�z�f�ZŔ�P`i��V����b���E�,Ҥ�L��~�/������|��g�G?�J��G��p\��ga��	�0������F|��+p`���ɩ�2#Ҹ�ڳr����6bf��w���x�3NXS1e���}�1>>���Q����΄f�P=��w���X�%�^����w�{�=ؾ}���g>Q��$�/o��uo�_h'��P��P�+�#b��=J[OLT&��rF���ÏJ�j�&FK�2�Gl���[7`�4�i&�T���P��麲���0���Bu����r�f���E�9���{����}���PP���y����r&�
l&dٷP^7��XU��]�"9(U�ʱ1�}�j����h����u�NMCHv����7O��㇓:�Ȳs>h����*��4:cŎFb�D�ן�BQ&'v����V�<��D��6���^s뵞u�3��]T�.SnS�wR���!:�Wf�n	�WL��J�)�359�YS��kHA��,��+V��_��(2j���EǷ�Y>wڲ�T^�6I�l�Ēv��s�*�LfU#o=�I%��n:5�a�W(��3f��ֳ�	L&�Qz�V]�'�RF6�H�|����̨�ʫ��
D��Q��_-*J��D��H�<�T�W$���]	A��� _^O����7r�e��l�6!p����y_�aB3�I��LT���UZE�������<2�ﳯ��e{�=gE=k%�>�9 �'�I>�����j���ڋ�������3ٯ�z����R�T�BH��8S2*?��Q�mɮ�^�
z6�^�l�XD��/��hO�$�[ߵ��~�D�##����֬�VzS	��� 1�	ɞ}&�1�R��p�@+�{���ǁ\Jq�𶷜��
��c7A�����4!V<����[]O�&1�q4%��b�;<#�6#7��y����m�� R��G[���v�ї��3�{�#�D�
�}������J^��H�9j<���� SW���z���K���6m�5$�T�v�g����?�RMz�	$�'�"gl�d|��p�k�3���!ȡ��I<m3	���AH2�N����h�ze_��>���j�������b?����{$��rHFGT��m��Ac5��`���bL�}2*�1��8e��Ҕ�7Pe���DciM��hT::f�t�j}��&��^�e�@sV�,z����h�L5�RB�#%-�~� .}d��SM����S�'m��Ǵ����
8��o����w`:7����ǿ|nڵ��!]y��]��v0�&��EM)�[T!�Hy�v���di�=�m��܃�7g�c×����ib~DW�������X^XR�ߛ��*��1-�`�� -"�+H��Ɍ����W��Vq��p�Ϯ�5�����9�p|�C���݁�!��}�?��J��S�\58v�Y�h~�|�፯x&&+�yE�`��Y��}��6�ݘ�I�e-�gu�hs�e��}HW-~�;�J���n���v;z�66m^����ux�˞��;rM{���S>u�*�Svblݔ*���� d�0�{�X]D���~� ��)|���a��Z���U\y�5��]����Z�i���#���#��:RQ�Ƈ����*��ꘛ[���*��~��O��C���y�#𥯜��;&U��%-�.�g�sf��ְ~r�rE�R� ԩ���M�.ϡ�8��Q1}F�\���e\��+p��<�'&�wL$��Qč�s��"�^�j����y�ڽ7������}�܇f}�6O�S��0�����F�����;���|-Le�)�Ŕ��G��z��(MR����,���23btfr�g&�m�$�ؾ[f�a��&F�A�{f��[�qF�V,������,���`����R����;�w?������\��6�v���!�;�K��eS�V�Q*��xO!��No߬�.�ۇ�ʪ���@kj���EJ��"�H+�f6�`7���J��U�RS>�8P��<1������'�\0�:��hODb�R(� ��B��F���P,��W�&��ae�)�)%24P�X��>��{���20�&&�hF����!U���E�=5`k�Ī�V�rӞ8��Ä���*p)�H�-�}��Cɉ$��H+�J[�H=cx��$wj�솼��E`R����6[��M2O�4"�'`�� ؚOe��o�K�b�ص�գHz��	�;�U"�&�<d	�*�(�������5UKG��'��u`�`zK]�"��Ś���sQ��W���xuëɶ�c��	%;N\{Sy����M�b̆L����J�{�}Q�i#��5,)�ˇ��C+)�yCI���m��LT��6�:�ː���	Q�����u���*�����K��fJ��.�ۙ�h��^݉>�H�MaDN�S\��O�f����R��[}��Q�������$��g���u�-@��4�Xa4�`%q�v[����y���|Uhm9�m�tԟ�V�zB��� \VI^k�c�]^�Ȥ���Fa�!Vo�"�,|O�ٚ�������[���`B6�y�<J�D��z��pi�Ϥ�TV��X#�B���>BlR4r#}vo�x}�ḁ�I��D�Z�*% ���U�c,Z��j?�w���?Q愨����gg*��0�6�dW���tgiW��<i�7"��#��Yؑl���}vվ���4�Rփ�*){<�C9�7E�g��܁fG�.s<+TI�3��vMYE�H��������o�!�[QޣVH���!�~�r�eu����H5dC>:���q�k5��j���p�bL�LU��vU-m��F���k)�x��}�b�UcI�=`�`J���v���UL��)���Gn�����I�5��������^��iW�j�J?F���&׵L�����r%O���4�9�7��0]>���Nz�����5z�w�3>{����x<��O��GlHX�Hҳ<�d�dS[�R��n�W���t�.�p�XX\D���Ǟx�zL{�6�\��,�q x��_��71G$�J"�5u������!�ᯞ��)K�ܔ���[����܊�Ŧ��A�A���B��A�l�W����l���laqi�.;]{ذa'��-x�_����U �_v3N9�KXi�1�q�n%��8
k� ��
�v:+4�ģ��/����	wݵ�>��t�]X]mi��̦<��N���>�Q��h��qv�ދ����n����%��,��m"�k�G�/��d�dy�c��*�ſ¿~�G�]�]0-W�JVzҩ�u{h=��h��ŖI��|^��G��g���,ᓟ:�_��
6�l�3��t<��Gbrr�R�n�s+���]����	��۷ľ��177�a��~����M��S?��=�(�����㗷7��o>�����ܞ)�-���H�#���#V���c����4���kE�c��yv6�M�㘙��H#E`��G���\��N�GtX�V��MP�?5s'�#��(5ͣ�bq��{8�kn�w޳�]U���*�R$Y5�y�a$���Vd/�m_渘	���bj}��)/�6�f�Ng�V�@g�aʆBe���9�^��:L���YAwC���-��zKK�5��s&GX(p��X��@��貇�%�n���^�Ϋ<�(륵{}�v[���g�^��(e�d�EUk��40�M�E���`���.���x�A � u�dO�` S�3�K�ȷ��V��@���2�H�L��D�{�4��l�I���&Q�q Z��SWZ��VXEj�ʽ9
�E�+2zO
�
�5��b�9�����+f�aU�i�sz^�l��z�%X��䖘D�h& œAJʳ�%�����w�Y���Z�p����>��2�Ej6�2�|�YE��p�^����m�'�>N*���3���v�<��#�^h�'�n�P����GsW�8o�c����ʸf�����8�$�׽��J�i!m�g�/V���V�-'��%���<���G3v�{,	j"���;����{����>x��IL���)��㽣Bh��OA~8�S�4q�N�n�,�W�׶�N� �t�h�|-fz�R�#Y�7[�3��l�)�I+�NM��^+qLV|\{2������艌�X�\�[1��S"��.�I�b�nTB�7:L��(��dM�6{Ʀ���y�n�y��hF�xC�cQ�U��~[9A$�u�f���]	O� 1��6�����}�m=L3yB������B�T��H�����؛L�@Ug��L��X�}������Τ��q,L��=ŦP�5���RZYvp�=��։�.ˉӳ��?����eA4�����"��z�]u�8�ۙ���_)��R	H�
�w�;p�
۫��7�?f.�\� ��x4m$(Ռ҂M����2�Y�8#��	+4%��S2�C�}�ͦf��.����j4i�����p\J���yF���@wZM��C��, 0�W��9��7b�Ay����{���r��^����g��5�c7Wq���;'�}ЇV�'����pxǃ+�����݋X͏�Ŋ�� $X�O�@9�:�����A��(�T	2�b�^����]@c�}�V����ǔi'��ӟ�Ϝ����x������58�荩<�?���Pi H�itș#�|����#|��c�\Ku�=���G��'?�/�{�3�L���O}	w�ji\m�k�� F����RÁ��b��y4����ӫoF�їA��g"�(��K��yP�GciT;�� �H����
�m���_�2���� 4`JW��݊|���+�޸�c�t�����:��:h7��l."�]���³O�4sxw��������oC�3��j]�t��mزm3*#rw��������=�m��M�
CT�9TJCw����ރ�'��C`a |�;�¿]�c�-qU�~rJ���0���q}u��=2iz�;�/y։��$�`~���>w���&,.6d 41>��;�`ffJclz�\�C��~�ao*��5���N��O^�1ہ�O~��G'��5��mM��[?�~q#�}Ά��\�|W>��$��VL��@%0m�Vbz]M���?
;J'G�~��*-e�%]�4u�q Y��D�!��V���CU�)+%C�#qT,�D�=�R����,������܋=��P���4
�����h�:(���Ǡ^.Y�t��2U�v`J��^�FV���^Y��_�S����8
���җ�����Fʀ�ά�7��r?��b��t;Z�]C���t��ӞeqH:��r �]�Q��Y����Ɛl�2��C�m�pь�J%�&����v��밓gr�6FT}:Y@@4�:,�TS��&����{��(���9��	�;̺���G�!z�`+���{z?O�<��j��Bj�U.�2 * %{ϭ�8A ��Ydr *Da1�>m���qKT�g<F�l=������9���	y�QS(�d���	P��9Ry�K�2,��X�jkɄ%����4�w��tfơ������Cz�jF���~~d~���7�L��B*i�W�-iMRC_G&Q���Q1��6�q;N�T��W�S`l�aP!�j�#��N@�y��I�R�C)�ӼyɌP�����lE)������Pz�RX�`^U�1F�Y�W�%��$=�@�������";�L.    IDAT�Z��G~�Ln�ޚ�;���	��VLS<I{6c�Y[����0��('�Ԟ��N�>Fcl�\�1$����,K���L�S��{;P�m�a�g�D�0�^��:gb��{6d͠�"���R�xa�FEQ=�]ڢ��Iߢn+Zun�T��+Xb���0imj>U��5<[�{�T�e4����9'�����O*�t_��p�����^ٙ��sˁ�+8�sb���${]����=�)�r�H`M�Z�)�F�_ό�J�rĤ�B�?��=7p�Q�0�LP�{�0֫��U/sP3$��H��3(Γ �����E�b�F����K��Ҋ?'b��V~��!��Zٔb4me�å&b>��"4*� )n X�R�I�z��4�h���mu�b��TFil�$�՚�ݸO����!��_j2^*��H�11Tqv��h"Ȋ�Z�L������9�iA`ʯs<&�9.&�]E���㷎�����1�� ��?��SϿ\R����9�:�Mbw�eQ����0����>��"����h��`����yg~;f�c��~��ci~/|Γ�Oox%�9iR�0~ *�FR�H�s{�8�߯��.���UU*��	0��ގ��݊�Ov��Ѿ!���s��,�ؓ7D�Z^1ɭ�/~*^�r�zȞd�;���z}��(SY�i��Ye�Z4�,UK��*)��S�3��:0mtG0�q'��Q��Kd�Nq��m,�Y_@����v��k瞢k��/J_�]�`Ϟ�h��h4[hw�(����sؠ��.�a��̣�A�����0:RE�\��H	[�NZ ���尿|��k𥋮��2o4{Lg�3��4KLz�X��w�ty��'����ɥ�x��ػw��m�uc��
]��;6p�X�y�Z���Mܛ@m�����߿TUW�Z��,m#�j�ĉG3�c2g�Ɉ��1g�3�HPT�@ ��4�f��m��x\5����"K�M7Mo�k-���˜k�����A�8�em}��<����u_�u�c8�G�׉����1�bwg+��.����a|��~8V�S���(z��J^�V�uA���=���^F���k�:Ϻ�x�3��g�t:N���� ��N�W0�jŨ���`�ܷ^�:��^�
|�"���C.b��9�t��ݞz�7�/#>��~|�����d�}� �� �=Yq%� �����U�nGn�;C�h1�S� 9(�0fU��^ܣ�:��^��q��v�F��ۓ�TUE��%I�7��RV�X�c�����w<|`���ם]g8��E�H�th˴(������X'��r��f:�|#��h���z#���;Do8�g�"A���-a��%���s��z/C��j��di4#� � b+�Lp��4׀d�d^]m�����N])˞U���P$F�J� �L jݩ�V'X� S��9iϊ�0_��j��cҷ�����!�Yٍ*��q9�*�!�G�~��4�Իi��?�9�$M(dnR�Ȇ�.������M�P�I����G�����Z�� ����c�<���Uh&�f��U�C�(#� @�h&��wIB�oY���W��t-���s���!$a
�=W���[zW[��d�����>Մ^�H'�%���I�di����e�ss�/�V+I?�!2,@2KZ%�ωWK=�ެ@��|SY���gY
��}![*{�'o���o���G���LRU�S��'Ūb�]�����cY..`+9wVM����$���1���D�SAY���{Z��B�IŎ��bԺ,ϮQ5�\���F�`�C�z�49~�4A*���35��!��\c�-I�8zۚG}�|�͸赠9�G�KB;��80{��/IB���:�̀�{����Şt�FkNX���tX�I�4���2��;C���'�ڛ��r�+�?1��ۥ�]~oB��h4i-T�/J�W2�qh~�k%e��J^'����u�*�l�$���3�E��=S�#�(����q�+�O���vetD�D�!��L���ܺ# Gc�e���Lb�^P�.W,�����َ�<=�z.�8��_a�[�����3�ˌ��DoW���0��~������]W���b�;
"˹�����[O8��ݍ7����̎
x՞��h����������Y1���a�s\m5�W`�����(a�,S8T��e ,x �10E�=��	Lo�r�������� n��mq�܅����U���k�}���y�
�r_ݟG���|$n��o��?�D�8`!c=�۞c���/��4d�*��>���T���"��hvB�=�1�Q��K��+�|ӋY}���Xi��١VIceO+�L����\�ڿL�x�����L\8��eW^í��RDy� ��!��O�X1}Ιa��ϼ�#n<�$�k1��Zõ�X�80�WUY��Y�>[r��v�#6�N#����o���������ر�f0%5dO�f���c9?������C����W��zJy��R����޼V�F�˒���8��^�Xg�}�j�{��B��W����1YtL�_ʤ��doLX0�n�0�����zg1���N7n��L<���kNƵW��c��裀���x�n'}�p���@ �\U� ���STL�<t�)V�snюɲ��_��yw���������y+�+UM;�!���o�]���cM`��;[��V���~$�ų���劬�zo���������ގ��p��溃����N�C}�X�=H���L�1�ۧ!�f1������B�tKá9�Ň�����G��RX_3��l�7҆$g<���^l��h:h������Sc=u�����a�;��{F��FʊA����"Ξ�Ħ#�?ASI�l�QXU�3����T\�|��C~�,�ʬ�H�I��zu[�+)7s���J�L��d��Y�.�����d���C$�`��<ݬ�e���U]����M�]%E �*Q���rz&�M��I�?/�d��{��@9ώ��2Iǁ�)A�.�s���R�	�X*�ؚ|n&/U���-y)��~����A�S��s��Lg4�+��(&�RV N).
@��=q��	,��B�&hb.�UQ�w�~[���>������˔����"���
�q�SV<�2R�=���{��4�$��:s�:���O�"j�k���AW�~����-�����B���X�_xf0�jm* �5��;�;��{�� �8.WFr2���0.P�g�`�kQ�)O��6{B�b�cB�1�8�VƓ�)�}���Sgo�O�fϻ��\#M��w��OW�D��<�5�mV��R֬ev���Nԓ.ҨѳYֈɎ��'0tAb�� �WqD���ݻi�Vǉ���S+���P3���l�����,�AdԀ����#��͵����ò
a�����Qh�¡��_�3�{F��	yGi1�T*�ّ��E���!cd�_;�h]��ź� Ő�?���U�t����<5UA8�EB&ɒ���' �]������]TIatԚ�	�,e�/b#�#�U�ҝ��lc�\'�ؗ�\g�4H�G �R��ZG�`6s�t?�ө�+����
4�kD��@�$I�Tsh�೉�@2��m3�l6e�~��Q� �"?ɵc���e�J�g	�/�?����_͢���p~1����g�6��%�&0��C��������c/ L�u����������.�$�� ҉	 CfS���;B`Ӌ�&:�s�g]���;�b�>�_�w�ox���p� �����g�������Ju�UVL �h�6�`ߓ�q 0������}k|��}6VL�㋟wC��_��z� 5���}6��_�ָ��%]yQ��񉙪��8v{��{_���g���q�N5?�����gR���aWիs�2��.j��{��������8~�JbY�k���,F%��lr!Z�s��3���߼�R^�"-t��R�������?h�>��ӥ�ű+��#�����/����)4��z���bi�/T�fcJ_c~>������~c|���̞��Ϝ�����L��.	�9��q���c���o��l�����XvN�tً>,�a
�7t[S���1��"Z�E�{�t�q|��j��}}|�Mg⪓;q�ɝ���á9�� ��'��k3��oN7"YLM0*�Pu��ܿb����5�̐��z1[G���8�������'|�"�VяvgH�W-U����F�^��4�z��G�u�}Q�� S���,f����I�b���=�oe���Ul	�t0Y��j,�_1��ɜ=�Ӌc�@�t�y��`GC�;*VR&�[\����q�� 6�K�^��6��+�IZ��{���0�R1��1�������d�,$��1|�pMG� �$@V���K��_P��3��>?�TRe�?ÿ���P&Y\�3��	f�<�1�3?{q�841K6���SNZ*;[�UiK�SI*h�#�������u�[;D; �3ˊ���YU)u��ȿ*M�������M�#�G��sH�@���?�T��٣C��*��V��L��S&H(��vJl������^�-E�;h+�ә�D����>F�Ve��,���a��J�9¼��W�D_�����H�L�h]տ/��@��'�D��]*%��:� ���fg��d9[��CH)��IV��FuN"�-Kj 0��d	ZsV�����قTc�H#|ߜM�î��8��$C�&(B�H�����k��-��KYa�)��j���:^��|��*��%HL1D-J0�z71����j���3�6G ��Zg4;Dީ�|�6B_l�3J5�@ۛ��Y�^+��b��%�A�(�h��T-B�r�t�NnC���	�Qs�&H��������~��g��>��E`�ϩ��5Ne���k>q�g���K��ۨ"��q�x�����n{s="���_�63[����B�����>ߧA�7k=�|}�q���[��*b�T�}��kS�l9��?����S���ߖ����p+xǠ-o�`��ߕĐ�-ls궢��-PjE��$߭8!{��<�b
�n�9_��� ��q�'c�F�[c8�.��(� ��k�{n
���@�8B���FM���=����#s6�@��x ��$u�v:�#�����x���x�,��I{��7��_�q͖�i����m��zl��|�s��_����ك8D�)z��$Jv)	ej�t���T��T�@�/� Ch����?{�̏�c��W���W`zq�w�F��-o������[������6eVK�F��y��ϣwf�{�O�����!]_щi��y7�k�eq�s�pt��������ɸ��M,��W� ���0�om�����G/�[q�]�R&#N���d��?�ELfCQ�@lV97�1���~���¯���q�57�"�� e�
H���M.r\�MW�g�5q�媘RJmp��܌q��<v<���H��������6�9��<t!�����[���8���؍�`�
H�&a�C�G��4��ą��o����+b-ЗH�85Ɓd��A�͊h&�$>�C��2ɋ����_�7^��;�=�*f�%��^��F(�w���.��ZF���|��\��}���g��O���;�~ )�w�����W����[�~��:��+*g��\��gV���p`���g��M+� ���;?w}���ȓ�1�é���:�[��PV�"{�춣���Q/� ���|����P}lGk����琢�٢���gw�[�6��mz�����m����h��X����cd�c	y��e�-�F �H[�����SH�U��>Ӥʌ2:�aXvDw���F0DB�W�W��&%�b��������!g`��Ǖ
.5W��2�Uәb�7[eTͲ� #�SZ�������A�E�>CKbiRSH0Iuhr�DWr�L&����ǕB��>�"�R ̱=b0��%N�����1X�ExmxWٯ��} ׿L�3�f��}�@�@�$��^�����Y��5��%|��2v%��;U�R"��q����<�r�|���*�JD��/Z�N�[��֞	��`�X��|{t/��d���9�ɋ@*�O0-��o󨸪��̙8&��d>�uV�2q�U.��sב�T���HӖ�(���=� �*����Gl��**xH���ҭ��3+�~Ӑ4�
��L��� B����`����7��8۸�	�и\_n�ު4�����f�%?�1�>�h�_xv�w�ɤ =�V�?qK�*�I5�C�DV�;��+�)�U��w�C��(����BI������6�f�!�s��@C>U�ʹ� � \�u��H	�ل	=�C�a^��$��7�2�ǒm Cz.G��Ŷ�j�
qy�I��,H}��>��ڣhD�w�u�"]�ljv��Kc�I���r,����)���w�쁥���:LN6]�KE:e��OY5UES�@L���H7���f� I����Do�/��\��X��PV�$CR|(�9�Os?��+�0�/�ι�Fb�Ire2|��È��*V0"J����_�Nt��vl��ݦ������������a�Q{�D�&��a,(��$�hSm�V(>�����B���4f��	�P��	�!3\�fl[��g�ߊvE���ZJO �Ŵ�g,[��q>�вZM�������O�������!�}�����������)d��>��IZB���\��\9�u:C.��s�٬b��d���ў>/�R���u�A�Yιo���o��������o���!N��Ԁ&:U�Y��X�4H�([$|�C���"~�?����$q�ج�Ͽ)^���/��tt-%0�������o�O?q0������R�v�)����Ͻ1N_�����e���|��᥯,A�9�q)!��CI��b���?O�K��;Xć�~(��阯��{��d�5�qHؖ�	弫����X;����~��/{n\u����{\�_v7�閿&s\��SBQ�aE|&��w �~߇�������O=��et���j9(�<�  ���<&��v�3�~��{���m�鼮��<l3u���Ɵ}���:�_ÿE(�>{.�?����w} z[WŪ��-�����M�;W���<�El�7q���8���g^Ϲ�ڸl�[�vzm��Q!e�v�����/�gM��[w�f��l��܍�{�M<������}*>pzv?�3 �~lڽhw��^1<0h�^����F.Z-�"�	�=��(N�:8�� �S�d��H:Я{�a�葀1 ӊ¬[v�u��	�����(B�;�U�ZTO�v����6+�K�Kʭd�"M��ꈿ��Q;:��3��	�8� L��Y}���`�+�P�eH"@b����y��ɹ��t�����W�E�8���># ST�JR��4W��2S-���zZ�cg����1'�i�$閫`ed�b�D'L�d;%x�j�QHW嬈�;�p�z'�'~|��č����"VTaUߨX^[�1��R�$`\C%�L���)=%�M@�f(Y��^4�x�٨e��Q�iXSyt�0V��8MGT?S</- ^$?��C�P�/�<��5Zyy��%��aZ\F�����$��d���bE��s�'�Q��0��M A�ǟ�dH���tWΪWh�;�E�Ѯ�"1D��քt��!OI��`�M|�G9��&.�NԙĩTh���h>���og�#����򹦫-�+ň�Y|rPoX��:?]zqٮ(��=��u7�J"�Y��?[�ۗ^�7cWQGx��~�	^P�縓�C��y͍���	��I�O����5ch�k�^a�5��+Į���1�0�Jv�$������)[|h6��>�����:"�6(�׹��N�lUO�?SZ��r������|3��OR��P����jt�${AR��3�<�$
�t�A9UB�Tr�wV;u	n��f�n��k�=�u�rs�[I�7�	���n/����P��#g����lȹ�)������֯Zt]RYpm�J͎	x� )]�z��仳e,' �W���z �9������n�p�f���RO ��
��>o��7    IDAT z	;8��0�c\�hWZ��9�f�ێ	TS�6��V^����ji�
u�rA@:�Lb��VaG#)؀eltR�i���:�_j����E��ؓ����c:����|*����W�?`��f��৞�7��o�=OLb���5�r��K�dF��1e0��s�+k�3�o��˘�?��?Z	L������/�����~�Wc4Ʒ~�߉�|�W�V�Q��������c�˿˭ip4�D��I���>~�=w�x��h�،�_xC��U��}��!ް���:^����'�0���v��/X�b�8�����lf1?�@�լ!��ITb��ޒ~����_��c�N�P���Rt���E��V���^�7�(c0ڥ\s�"6��X��l���j9��t/��sq��q�5�㺫O���Ʊ���p�m��傹��F���s�Z���BPs�����h�/Y���x�����<{�v�ND�; ;�uc��ܫ��ii��<�����oO��ϸ<��7ƍ�]W^~"�����a�>M����������a�:s<I͢���q�pO����>�{���ԅU�����`��:�0�I��{{D.�b�<$(��4N���]�<�x�W���O�V��^+F�~l��P�h�����~�5�o�|����Y̖��-1u��ӈ{|"��}$>����ӈ�vDW?Z ?�5��Gİ1�ƪ��؉���G�X�}]����la��d��<� ynh�GE[�È>���\����LPǣ�L���1 ��l�T���>zN���@�C�S�+����koT����Tʭw���d���~Yg\U�>V,�,�W��mQ*	*Ա�O�E������r�*(�
S4$"�~fu� r��*<��B�=u��e�R��	��`xe��L`jḘ�ԢvI�l�5K�3�Z�ľ+7KX=X���9Kʉ2�`U�{���{>0�Gq��H�a=p��ERLe��}6���T�8"%�f���-���J֧?��R�;������d�hY&�=�4
C�
7���U�$�0?K�P�F	Z;�r��mJ�t��I1�E���܋pU�^��L�U����j2��Q��J�"�1z>�
*� zW��^j"��=� &@ٿhRHȰ@F"m����P{@���~��8�*U���ْ�����}����T�W&V�d|�e&��;�iW:U��8�E��x����J]c������2!�ʧV�kD���e���:mEH�R��zM ����11/�Y�g�s|G������Ϫ�"�8(TtL����)��h�&b�j4)"��� ���n��^~T �'V�_�NJY�t2�ʽ����HA����k.5"Kє��'IDS�3��kU�W�~�ٺoIԀ6 �G��o嫒#�¿�S)nP8�^x�>ù���Ң�P�*�3d�Y1���Wf��H�8(!��b'U:>�9J�c �oGfy�V,�J��A��'���`�%���t��{�E�1(�>���%���`=4��h��RG�nV���PIO���v�4X�:�/�Q���3�ͱ0]�3��"�����<�80�r�:����^(���|8�b
���V2v⺥0CeV�z�qk`ʅf�F	4�C[�
�t[ˋq�M�ŏ�7Ǖ�^��j~��f�����	L�{z��(f������@W�R1�܎S��q�����)�ެb��d\�+�����o~M\{��ꃃ��/��ߏ���;����7���7�O_�[��+�xnXk>;�g9�1�i�>v1~���w}�8/b>ݏ�b?^��g�+^�O��^�>2�O<���������ڱ7�P8���^�v��e,������z1�}�	�T�SlL3����~ ������.��6X���%$�z�!
�JɄg��I4�'O�'ߋ����:�3� <G7�@mC��c C����2�_Q�4�Pu%7?��d�pm��(60�Z����ҏv��V��S�(�_=
b�8�t~�9F��b�<`�i���~wC�t�sMQ�C�'LXS����E9�%o�s�YCF����7����u̖ �;�naG�Z*�-��)سLK	�2:�I�;���-��S;q�M��sn:7��"N_uYtc�A7v�G49b��iT� �@����,�*�!�=[�c2[���,�z�����'�d��g����y/��!4z��w�`�o�f��6�X�PIYUt��Yw�"F��)�a�ίE��T�����	��~��Ħ�2'0E�<�q1��pH��7��2��A��{4!� ��ڨ�l�e:	A!��'�S�F1�KIȚ�e�pRt��I�Ad���t!�|OB*J>S֕O�u'1Y<�D7+�d��I`sM�a�c_�>(��u����j�V��'�>�L�%���� �
R�փ,c2և��t�+P�2��2�ԝ�V�Y����g�R����Y�Q�V *]]5���A�Z1�u��ӔZ�ǭb0�%���j;�0�|�ѣ����U	i޳��t�ĳ�h&��"�R��,�婌ͨدj L��,���Q�(�q��ܬ�hO4����q� ��������%��7@��g�"^d�k�k3���K��2:U��>Ҽ�
�B~XF��Au�ɿ�)Af_�_��"�L(��<�"��PV��<�dA[E�g�$�Πz�� I5U9�������Ji<�f,��~��ڤ�#�)�#�~/9lJ�+qΦ�j/6�V.�R�$aղ�mC]V�%cO�Ь�Ir�
��v,��j'H���L�?��4�$���8��R�0�tu��+g�][�O�W��5��2���Z0٫�D[��*��j_'&p���p�t0��[́ҕ���e=�ŭ��H�[����)��\0>�ed/���(Ddk�*�ճ �ؑ03`MJ��z����[	���ڃ���a�Ub�ds}����������s��:S�lk1��Q	|�@���?0FFG�ؠ-kw�������ƹ&C�1�O�h:� �@.�X�r<���z?��������$FvK���x&����P�Av�&T����W�T�� e���<��i��s��5�Y�Z�0	@F@����y�%�Jf�0]�����~��L�l6��G�o�����<&m��Q�B��<
J���!���)�� S-�d� ��? �{g�K�{]���e\wj�}���c�+��}��o|{��O�k���_��~U\s�q�xDR��^.6-XJf���{ p]>TT���e\<X�G>����O��=��U\8�x\x��x�-���_���[������M+>yv/����ӏG��:`uz T]�HL�,�R�;�g�$1fNv��'��^iaT�4�\]���$O�e����u(���i��GV�~��g������V,f㘍�l�^�Z0 RΰX�R���a1x�\��	)G��a�w�D�U��> ��^�B/Z�B�jn)�#�H���Ă��K�:�:`��1_LY��-�7��A"�חϞCU����Ըg��+*�A�<����{๡b#q` �=l�������A�Z���ɜ:X��Wщ����iߎ�������DPz�����Q�z�����Ҵ=.�H�������i�7>��r����MǋV\���3�^�����?�d<��A�6����X]�Z��P�n��A�R�U@����A�Ai���ml�Η��r��)�E ���Cu��Q�� ��0i"85��_���9�#HN��aZ4���pk|+0J#d(��!O�S�N��\!Pᚄ#�Z��P^���
#'�"���� Wӈ�1~�$
F��t�*�iƮ�f�¯"	RRP����`Ꚇ4���eHz�g���!̽��z�q��L&Jr�d�re��_Ӹ"�ݓ�F�e�ټ<�m���`e��z�zfHXEe@�	�֗
OJ&��+��9��'�ʽ+0�g��5�&�$�\�uҌ �J~%$��Z�gXd�M����g3�A��~e��T��5]R ��	h���z@Nu��x$��4�43��g6��L�]��[Β�aV�1��K~��|Ou�F>�b0c�U$M��oB���U[Y��,�?��yV$�+��;V�@`�g�Q1!�5�O0Zg�W�%э~IV-pp���i�R��� ����XP���C�lJ��6VN�.˧����z|	�D�⇠43M]����2���}�)aN�W�fLZ�u���HƵoj�m�R�����H���ŔBz4?�����_� ��.��v,}��ڗ����_�Q��r�b��g+� h�J��D��I���� UaP[z���ʊy����|�M��fo��,P0V��)��Y�.&ei��睕W���zC�F��d֫9�����N�/�D)g� ���6Uzv��?#�b�� �R�bb�%=f� ��ڦ�wIp����3	by�E}!�r�E{F�z�Ck ��q����m��SNT�^s�W��7:�؊G��:��t*���ԆD����t�1}Xyb��Z��6��)3͛8-�]|�< �x7+� B��>��.��]�����	"�h�}�#�r\�t����G�Յx��'�Ǿ������>o|������1mo��4�<�U���sT5��UUT���&-�L�Ņ�����x�����k��˷�/�r����w�a��_�t<z�|�<�W\v�2�>��!����UZ|+U QɄ��?D�Hj7�3��8��c2�C�n~|p.�?�`<�c�W}w��/��P��"^��o��]�����b�
����)^�b6���l4����6��m�Nd�DC�⣚׬]�Å������If�r#"@�����$��
9*�q������Z��� }�B�t�c˄2	�Ò|>*�Y���*�.@"]��X
�7�E9{$k&�.�ߊ���2�:�
�������-�t�3;ToW����*�����BV��`�/������#��v��G�<�Y�ݶ,�HxM ȋv1�-��x�3N�-7_�]s2v�{q|g'v�bw{HPZ�F���盱�/�k�e���&�aP�w���i��ić�~(�����s6�a��[��O�[�o�3���v �[�՚��(ɀ����'�B�m���D F~�:��~���瀟��'p��>cI�� �I���� �3�f�'����|EL �;��9J�Ny��R�j:ULq\�ʾ�;��[��9�<�ȣ����X�8�	����69�ק���({�m6�L:x��5UI�@ެl��*���)�n�XAyY��+qJP�$�M�&ǫRa�'���'L��s�C.c��"I;>���V	\������⨪%^��[L<t&���5�{ӡZ䥍J�H��\LTD��&s$ni���@O��3����S�4�Le�-��r�<KM��U� 8��g���Β�Fk�$��,q�������jd�"�Y�����3�+�gz�+�')�,O>+T8�Ե|}���B(N<G�������v�����c��srmy�5�"�'�g��I卾�9GkC�J�Di��M�/e�b$7��MEϴ�P�Ğ������p�� ǭ�kr��|r�I�(�EQ@����a��"@o��Uk��g^�5칂�l��.��Ha**|�/;�By
�T�y�$e��+��q�݌����v��_�=��%`a5��T�0SH<^\%����l��+,��<�+]�����8��G�T/��9Z+����y�GI�l�p {�ࡐ�RE�b�o�1�~�"	�zPd�	Nk���.å
X"l~b�מI��WG$#�����-`�@���NU�t~��!��=�V��@!+N*2�{ڌJU?���ޑ;p��c�Ñ�9K_j/��&\���I�+��J!��Dg��5��!�w�KL�P%E�2� ��J����|�t~.g��_fG蓝�
?�Ɂb�{�C_�R���y���1�B#��JR~��g�Ƈ�"���[�	L��Y�Ǐ~�KLQ��3��ζ�����1�l�	dqIE@qF��;��*A�?s��_�15��r�X���<��j�l|ɭ���b\�;�P���sL�W������ �~����U�,^خ��wӶ�A`���
�`��*�
��5���|\f7^�ï������L�'"^� ��8\���}T]��W_Rqv�ԭNflV��Ԓ���J�6TVM�د�	P*0!Ub��k���
3�`r���N|)�p2�썂�&N��C�3Aҁ�E��wgsj�u�VÌ"9��04qV�?=N�P�
�l�i>Akpɩ �#p.�+֜��||m���A�}>o.k� O !�Z.brpX�)�	W� ����:�Ҝ80��̸NYm�Z���[�d����y�S悤	(�6���3X��0�S�x�s�����&N_q"vw�qbwDP:�l+qV��H�JZS���޽�?Q���faxoxG0�8E�鹃U������?�H���1V�0�=��<E��7�l�%Wpd��jZS�]'v���cH���N��a�3�#�-����=Ć �s9wLk0��4¡��;D��~-'PL^��ڋ?} ��
'��s�
�Gʤ�*ߑ�c9�˧��ˮ�A�����}i�a��5�I-�F",F�VL�P	6lds$�̊oCN���E!<e�5�O���c	1�B�w�1o%@u�� �A-��@�&���<�f�x�:�e�$LkI�2A<��@ޔ��QW���˧�Ě�h��:�=Zu?��m�[�����&rB���dK_��7�	3���T�����H$��!�M+I���fT$��l\=�{�X(��zSY���B\O�mN����v͌U�3�RC�T?��kU�|Vd��}�6к�b�%�����O�C)=��0��\�ȄFs�1�Hꙟ�j��J�J��g�f�tϹʻ>�ϻVq�|�@\2�<j&cN��T��GHf�7k���K�w�着���#.������C���Y���@���_z�p�d����`	LDHP^h��E%���eu�.I6�T?��R�S���})�"�nT*�:R_��U�Z�]�Ԩm	̥��x_@\����s����a$.@���~J�Q���N�m�x�)�Z�K9�M����@\���4@cZV��s���Z�&�ݗ/��VNx; c�c�]�)'w�W3S�N����H�M�����\5���j#�,�$��sJ}��%l��s��u0^g՛�sG�#]�}��_,<�Ā��D�-�h�,@,��<|捲�yJ�5*ō6Ȣ ��Q����t���b|��)3��|w��Y�%���ޣrt�ʋ�Ȼ5r��H$�� H� [,y���n�3�Ji�Ɛ���Wx���x�Ԣ$L���X�t�Fc#�/̣�:������g_?���������1����?��ǀ��Zs��m01
}��K�%�/���tzp!��x0V{g�����|-���`�����x��_�D<�c�@O㒋�A�+��B�nU�6��$��!u���{��A6��z=���b\w�X���@|��|)����'������U�O{��(�ĜDS��t�e2�"���:(�e�Q���^���뛳��,�R_š���<eલ7m>w��1�� #7+�^[2�v�3�`����x�)@)zK�>.eT��/�)�c2��E䆪�5)`"D�3�i`Ev�	B�J����PR�^2Z�_,X�b�~�,R^HB0G�U]2�|�J�p͜=�6�nf�f�,��
��0[
@���=�ۍ�ۭ������[n�k�:'vq|w�.ۥ��W�#қL%���\ӭRc��0S�Z�z�g'�>}�����w �{�XoF��؟���k�37��!9G%�ߧ$��$F;z�F�Rs���!{F��X��p�錕Th�(Vu��8!�w���!��Ň��,�/� =�LY=���� gm|�ӭhooŲ��F}5�H�US�.�֔'gӬL��;p�j��)�С$ʤRV����%%��P0��>���͕���P���5C��~�H��'�P    IDAT���E:���$X}8	l���ѳ	� 4�K�"��YO���hIU�9��8V�ɱ<��6���5̅RnʯK6��T���)C�D/�Q&�$��S_���l,;,ra%�`�)���
�@dp�"�u/��>�S�A@�)�ʞ�,j������}�����4�1pR�?�I��R��}U\?#2�q�d���xgr�\V�\�g[��#?����	�{��HR��V��YaД3�2T{��b�����57�Vf��L7�ZV���b#����<��D������n����}���2�����ɘ�,\ULQ�]�-�:����[���f�x|�z��P&h ����먐s�d��4�z��f�*:�D���j�C}Y�lV�^��Tm���u�9J$�2U%)��I����|JD�ߏ�/�d瑒NMr�i�I0�W}�Jv�{�!f�dH1Bd��m9��.�f�0�y�H�e�� �I�VQb[u�.�$��ú�nʪj����5����R�Z�}\�OGv��M��T2uʳ�8N�K���,�u�A
Y��}*�RZ�+�x��{��?�5������q{b���H�;П+�~��r�*�I�22$��LE�h�#�B�f���/ ?A#��f`ډ�`�J�$�{��9�Ϣ5�|w{���%��P"�{"���9��`�4$uh����(�&g��y���>�VG���m�3jai
*"�ʚ]���o�Q���3�"�=�h�¸�Il�.Ɨ<�T��w����6��z��W��~��ƛ~�S����tbh�r3Z:����@�rS%&Y#S� �aH��Wqp��������L��O`\��)�	����x�k�u�������SnFھ����� Z2M 1��:`�ء57�Z\��"A�Nb���� n��T��5�����/cU��ﾧ6�zS���*�g�����'���h&5������M�61����y�6����"��\K��d6���Mg�n��d��@-�4��UJ���gs���qw�jl��� ��^t��X�^j�Ȧ�Մ� 8�`�%%
��,�N��H��8
VXPN��;kVTG�y� �P�����#72"���:�`��	 ��g���b�vb�ܘ�TU0Ɍ-}d��3�ZbB%v"�O��qĤ[}� c�k���f��v\�ݎS�{q����>�Ƹ��n���8�;��O��i?�̶��\�Y�2��l`������@����l�M<}��?��|���T����a�P�W��L���u���A�ҏv#��E��c�X�T�� b�l*�e�&��7�D����KF�t4`�)	�Ne�"��Ϗ�k�A��U,�|��M:d1����(��(֝>��8�d�8g��*U��>�J��rr���r�v*ਫ5�=�
�������z�d$I.V��\_̓�@�ġ�N2qf,�ۦ4�I�E�=I0�!�R��)�k�P��MgJ%�5���`Y��g�H�E��U?É��HӃH�`1�L4�D�6\o�E���d�x87>
�vIJ�d����0����A�0�I\V���\���gB�U�z�^6��&a�v��َ�Npk��Ia�"��,+��r��	9���%յ,y'���Ux%�������z̿Ӹ���*hV#�{��3����$	տ;*̌�ɠ�I�'W�k�Y`�I4�0�����,��u�T�{>����Y�*_��C?%-&��Y�]�J�����G �2�R94R�f�%�OU�c �*,�m��&l��s�eŚ1!s$�͵hp!R��]H�j�� �����d���k.��kD�� 0㨀��5��J_�I�l�!f:2N%��ͼNUu��(w��E� �?wu�c(�P�J���y�A��&�Vbo���v�RL"�g��k8*���J���gr��k�yM�$��;��XU�R�3���hr;�
Ќ�J�r�gC����iX���e�Uފr�� �@-Ğb�گT���LuA}�Ib�n�Jl}����YvK�av���w-��7�x��3Hm.y2(FH�@
�T]�}@�B~�������5yUowD?�ѺP�!���ߊ5:k�
�G��b�6�����Ӂ�����ۏ�;{4�<�oZv1�b%��0��9�Kb��U��݊�W�Ib[��x�M�ŏ|��iJy�ĄF�B`z��������Y�1Ǵ��W�J҅�S��@J��T�$M�}6����=E���ӏ���YVL���3�soyu�H�ZO����;��3�DND�͔R���\��Л��h���`�A4>�E�2��
�����ӧ��_��q����N�W�����xٿxS���"���F�}H-��jU��d��CT+��K5HШÒ��d��t
�&������)o�hr;q�D_))/�>+Nh̬��*����{1�wV�H���c�er�'i�ΤF2�x�R������ڨ��^phS�<�|��3$G�nm���YP�+��/�S�PZ�*�e8Z# ��K	�L����d�����
��5e�RU� �+E�*�`Q)�;�<�ow��c����0n��t<��k���(��8q|;N^v,�=7�7nc_����L9H�u��x�M��"�F��|8���?�'��Gwt".�t2���×!��l�M��%3С�1�k�"!���^����d0�e˃��.�RQ�����ܮ�P���4�3�L,���DHh%А��x��LF`wv�����PN� 0�g�
`�P�!z+����H�oĹ���J��j�@
�cr��~V��_}��O	YM���jG�?��_���d�}ا8X���L��xgՊI^��!M�T'�����
 A�T��8��Zd�q�0��Km� A�#�L���"�՘���O�>K��hNR�=>%��=w����Y��{eu�� &�F��%{K�ڥW��	�%��ZJW���N�������Vi��*��q�����!@`s8T�3)ۭk%�_�h>�T�+��;�$����-1&}2��>�&SڙC]jE�]z�J���1��jޓ�웆�9���u���٠�a|�2�"��
��|��Bp�de(׿��k�O�+%��2]�M^c�2�g4v8M��-�K��r��sMJ���/ �g����� E{��h��Y�&��������y �����*�B�K[���ZK97�W&��{����=Pq^Q�3�A��A�����~�Z4Yb���f���&E	�]=MR?S:��I-2�)����kƹ<D�ẓ�?�uU�$P�yr�ϴA��j(:�M��s��]�)���%vg5��W�����3V��KB/�G�a&~��]9΂	=4�pJ�C�fdf��E�&�W�M\��P���	u06P�zƎ$��(mE�������A�}�mTJћ9���F,��'�cL�#�R�1Wn�s�Y�3"�Hi J9۝&�SVJي���PG�̯QD �F��YH�6&U$�� �lo��,��K�/U��W��g���8\^��t"~���W5zL?'0Ÿ�|��x�/����0������t\"�B�����8��|��8�x���檎���S����c�1�_|s��Ǿ���#y�"I֌�T��RU����ِ�O��hM*lL�q>�L��\�l�߃˔\� L���[���`
va�~?���P����Õ-�rhu���*���%�6!*�<�m�v-`3�)���+����,��J�J� i ���8�c0�<�~��F3����X����%����C=�"Y- �)̼e��8",[s�N*)\7t�p~EE����H?mD6p�$�TΠp$Wp"uR�L��Qi>��.�� �.��u���B�	{x���A������1�.��V+�<1�3W�rD�3�q:Nlcwԏ�Ƕ���������jU-J�L���8��c�h������?��{��.Dgp<6�gK{�u��({A�����E�?� �){t�,3��e�X�0���f2���~t�s:��{�xC$��+�  hS.�	L��1���]�=��e]Og1�������ڜ��َ��V�� k���!T���K,����� sH��*�&��R�D��K��r'�h�����K��<���1��F�Cu"�,���t*5,�b�qr�d#A��f�ق�&����O��
ܝ"�3��3&�;��bXVH�%٧��dν���U�o�/Y���%4�ι��ɔY������)_�|~�ˍk� ���LJD�Қ}��@�Tܷ��I���]���2�Ҋ��_>W~�̉��:=Ɣ>:��lV�ӝ���,S�K�ّ|ũY��_h�Хe58M��gJ��_�$�%���d��?���e�Sx�k���b�Vi%]L��~�LM�3@��1�	m�s�ʷ�;;��~��o���|ͤ[�@����>�e��I�|�^�2�rf��$`;#{?1j#�h�<��T���;ʹ}�>��2�=R������p�pk�r|N�ʩ��A1�G_�vL�qE���!_��'?��F�r��ű��=�֬�_�Px/�ѫM����e&��b�J�z��E;�E��˳��FU�U�J%L�WI��P�O�������j�E�S*�T#�
$z���$5���1EB��c:�g��ǅ%�~^��&A�XE��K�gM�Y���Y~�=�>���5�U{%��e����o���&�?�9(�H��@"�mjlR�*+�T��5\G7��'��s�V�鄅 ������E�ٷ�Z�rU�"���!�q���A£}�&G4:��X����?s(I��g,�9� V  E�L��>iD���� �Py���׬g��Lc��_|�q��b�!����ѧ������[�xW��Ĥ STE�i>�:���)�|��T�9xXL.�;oS�/,�W���X<��'�o������#1��M�YZ/D�[M2L�@x��r�x4�#�O��?��"	�/9��b�������-q���؛���E�۳����	�fvs��˄���h�$IE>&�E�m�r w��X0�劶)2Lo�v�3�t�L�'�46��������mm�t'е�,��O����w̄Ύ��Ȯ��V�!�c�q�S��L�΍AP�J��˔6�����|8��������kL	VT��K�4J��d�:���N_=���0{VDT�� �]�^q?�@[���۝�e�����ګ�_�����ӱ;�ű�a��bi��>%`��7���_��ٍ?B�%�$��0�-c�j�t5�{?s>����~��Xl�t*nu4��A�̑@�b@@��-�!�r�F�p�c�������R��N���4��Il���p�d��-�k\��u��sϫ��L4>���g_����88��l�y����������h��X��z�H�`�0�Ҕ�Ns��%q)T����Ճ<�4��&B��N�2��d�����ُ��=��g�(b"�D���h�9R9�^%�4�~f�(a���Ia�S�tT`j�Y�(<#�3��\����s�҆N�Pk]��W�Vf��bPMNj��&`GR~7/}�j�Q2��n7@n&�>L2irU�n��V�)@]��j����f�2�i�{%IJ�� pF��1��/o&Y��p�~T��*�3?�bd��wia������ݧظZ<�@$!ݯ_	0Kk]Ib7�)7WB�5�^4m��#��z>\���6�����q��%W��ﳚ[��&5���`��h��B3����/�T�#îtMX٬�k/;ry�n�<?����S��)Oh&�yn��o���{,�S%�'v��)�x�"=[���һ�k"�g�a�q��Sr��	�o{Q��3/���\��N�S��I��w2U���7�T��(d������;��T�+��3U���_��������3�j6�f����ȵ{���y઺a���:��D��T0ZE�?��P=�i��o���ψ��K����|�y�c����,�d~^�=l.e�s����[*��ܼ���a�����
��dE>�Ph�&� p�5����'��Z�n'j3��B����oK��o	)�j�����3���b>��O��U�;�bf�R��:ɽǽe�֒�E7����# ��ol��<�	}��B��U�,.�k&>Q���%�k|����s\'�)�!��bК�p~>^pñx�˿)�Ʒ60=*̯і��λU1�ԓ�8����S�t4��b�[(I�\T��5��Y��\x=갊�"f�c9>��S�u_u[��e�0��E����8�	ց���,����[2,Q3.��)�q�l��3)�`��*���*�?����#�؟��;���=X9��b����U;h�3���@R��5zt�G����lqj�!4��.{�rQH����J���O��E�b=>�7ЬW�^'�iL�3
�b�DF���Le�k�K����`@�yFF�(��"�r�0�K/~n��1�q��3����&nHP5�"6$���c.[�A�A�f�S���a���Y3�5����.�0�B�3�YL��^Ĩ��;��x/n8}Y����	LOl�ı�����R`��fzi������f�`z�`ʪ��G�7yr��[Hwރ)�N�stI�����ÔR{0o�)A��è�&��Ѩ%<�X�b��
N6)͞-��9��i �����>�0*�`� ��c��f:�#l�q�ȫ�� ���c5>�� ������t����� s��@h�Sr;�e���`�9J��&淂"�����&���3ٳ�D�/5a��wW��껖4J���⊜�I�V{�gQd�U�{|��[�����'�d�6����7�	�Vm�f�:/��i�Y]�f2��<��=���3���$�ԝbDVY��t0�v�	�7�3R�Wf=��^�x���P�cL ������=��r$Q���Bl����#VR^����w�>�#��Z�)k�Q�7,���vW�t&D^U~�~�	����O����61S�l�'���9a�P�WJ��jl�VJv9����:$�V�U��`�&ǣ��B�*����Z�K�U�a�ߧ֟w���7d�_2���_:�@��j���X%�XX?z\�ڣ�Akᨳ��$���|&ɚ�i�J� ��fE^�����*�]�A�4�S���3�+Ζ��7{�����u�\1[��������7��$At�UYp|y�����B���?۳L+��E6��g��:6�3���������HZ1�{R��+.�u�LSn�φ"@��M�I�I��ȯM�
c�eĹg�(�<s�����s���WW�Q�� +H���s�k3��l�Vk���@הּ�$�F5�1��,R���"GOU�������݌%4�k���}(��]�RTK��'3��9�������-�AA^˞Ub�nd<ɾ�mc� �4 Ť�j�����|x�u s��Rr�������׃7
C�̑ϕP���m���TE�c1�F?f�Ͽn7~���%���<�� ��x$~�wǽOLb�I�˞N%@	LY9KYg0l:3����/%ʦ,f�n��	8N��ў=/���Ŀ���uJ3,g��!%�J%��/��876�H���H23� ��kA�ސ"X3mE|���G<��i'�ǎ1�Js���a4��r��,�p��B����|��&��c1_b� ����q���:�ڡt��� �`�*s�C/sђL�Z1o�j�ډN�#H�`�c�{D�t����wE�m��2��)˹�rT0P�G�@a�R��@7{o2�H 	�|8oL�p�frl6��͖���#;�����/KYrc�<��4����̓lD��G���;Iܨ�D��{4���k#d����5Xэ�Ϝ�/x��q㙫������頏$4�j��\��n�TmG�S���,:��� �8���z��w?��ź�\�B��a)����i�K$Wp��<��%�@)H�kN&��1�t���l1�q�H��@֋w�Y������	L�㹪�[ãux��m���@c�%��=��C�D�Gb0������06�s
@�?�Ĭv�`P*�)%�>vAF1�cVu�S�� %�w)��&&�st5�W�$��q�    IDATI r�!���ɪgf�&"�(Rk���5{;s\@�])���	)����-�e�$�$Ӹ�v���d�'�����M�Kl���Xd)�_�����b&"�
�]�Jr����1���G��U���1U+�@��d�S���gO�͚��4���1�%����z�$��6��/�����1���� ����+K�S�n}�r_�JJ���J	���1��%�C�AFy�&JD�MO*qP{���h�� �|��T%Թ�i�ǵ��F"��C���C
��/>�qg�uU�)�`G��

� ����x!K���e&/>�k�,"�[vd�T����G��$qmA�>��ߠr�|�}�$��M���k�4�[����������,��*V���>��"�}*��~_�/ŻB�\��aˣ�`5zJ�Y*m<�`Hb����V��S�\�����s(��R��8��G��!	�+\etIf��S������9�2��Y��|���Au*��M��,r�k�G�>��1���c���}P��������R7��w�AU$���J�B 	����W�lV9�&�m��}n����<g�y����ˮ�� �������lM��>��m6�+m�R��������
2 �.z>�C��J)s�m�1��8�HCi�����6d�)F���-P����5I���1��ȱ^�#��=�y��V�zvkoz��q\\(���w�Ņx�������R^���n��E`z���_����iL�#VL�h�>H����g&v��#�lJ����r�)�ep�D{yȊ�7��7���q�$�JsL)�+~b�-��v���'Y��C�c�m4��|kԧ
-lz#�8(M7r�,^�ē��؟�b��eES�  �c5?��f/|�M�w_�_ŵW��g�-֐�F���G����'���O�[F�3��b5��v�q�W�s�s=���=�~����a6�gV_�Q��g�#)��j�Q(0�2���d0![[;�C�s�b�p?��	7�|<��P�݉aw�������D���n�W���1�M����v7F�C5E�-�$���6���b��!Y�#����5���(:L�a
�1<��77�s1�Q�@��5@>�� z}����U':�~�9Q+m.H����w%�i�׋�pDc�AH�3*�ҋ (@׿��]��+��Sl-'�_��_R�{��~<�����g� `���ߍ��>��ا�U�?wk�����a���q~���h�G��^�;��[�sW\8��.�#f�r��b
$HW)�D��d"�XBj2ڊ.fp�Q�E�H��VmpV�"Z�M�PyĘ(HQ���rΗ��N{t�E(撒a�a+�"��y��Sr�^�	��~PT��X�	o.)>\�:�Q��wsT�W�n ~��f����9��#�������H.B	���M�����!CoT�%Ъ:V�`��Zbc�״�]��?RƔ���� )�iY��i���P+7��!-̞�T����uU�J�;�w�W�~f���f��Z:dܐ���EH$�����ׄ��zp��DDDeי� �Q�a"�R����0^�80ݻ���	�\S���6g_6�ub��^�<&Gfu@���D@����e�?/�ye���D
hP�`�+�:+(��%���^7Kۋ���˾��۽
�#���2�5��_~�ʪ�����B���DM6�Br&c��T7�0@:-�$Ak&�E����D�	�T�+rw�&�I�7�R��~5)O������e�X�0T֨*eV��b������h<Ϧt��$����=gY!I�k�hG[�8��#��Q��
��]��n�ɪ^���O��_�h�U^?�d�/����Y�T��� �Rk^9���)��Ꭻ�b-����"�?���u~�G�tI�5y�|1YEueS����p#5��&h_j��򌲤>�LU�?U��}���1)q��_5['�k��\��ɜbP@9�=��h��K2"c�HE�s��$��A�,�MԑO�������r?zq	..�]ُ���&?�9N% �� I\u��r�!�X�����0A»AO�lɱ�ȕ�o.��\B^K�������k��g���>Ap��0%jQ����8��2��o�����=~6@)c�Ϸ$��@�u1N�[���?��@!ڌ"��~�ܨx��<99��b���x��x�+�=��|����x���SONb�ފ%F&0)����5��&0-�'ͮ��h�y.���N�0ۦ���|��m��_��=��8�5�ݝ-���/�� �K����@&Jv���6Ɣ�,��� ��VN��X�/�>����!~NHY@ָ�w�����s��Z1؂$��o J�XM���V������1���*��籩[���;��]����b:��lzW������������8q<b@�g{���������Ek��?<���&�⽲z�q(�C�~�t4� ,�1<h��A��5 �$:H�f�h�0RiǏ_�.@Z7�辦�F	2�5��ۙ���Bt�J���n����wT����`�=%'4ΡL ~M��p{��KQ��9�T�`��8���p_��V+��[1��8n���.fl�z�����^���0�s���t0�b�[;��� ���;��i鲠?��(b`m����,ګIl�qr�W]6����"n}΍�k��ˏ���ݭ���Sy��W"��T��J�*��� �g�����h��to����w��O����X���TIq�**��ʕY��UXs�![;4-B�錕���r_M%W�W
�=|�tF��Ƙ���6	G����P�Nt�R�H�,���%or�]�&Z�ݏ'�<S����.t ��X�ŋ�!�Q�u�m�J�&�Wjp��Vu�d2��K^[��:��ZS�^@����$�T1�5�D�xQPs"rs͊��A�2�m�I��\�R��y+��z7%|iH��2�Ȗ[��Ϫ�g��J��|'E���R�~�lӽ
@��<���7̚ie"��G�P�B�;C�sG�F	�@�l��]`�
@^�-U�96��s��b�,�%}�I�.*	  ƈ��1��Q #L�\��lfU��ޘU�*i�z�O\�w"�h�fP��w")S�
�<#ЮȌ��dt���PX�ʾ+��2�MP���H�y��2�j�l� 9S��e��M���eT���U�4��=@ј���ѐ�g5?�<ϸ&L̈4��<п�=��3<csΪ*�gX�*d�dzP����n�HH���q�V�s����c��_Dĸ����l ��;�0RaQ*�Ҹϰ6P���lO���t0e�ZM���_�����e�$�"2,[������xyåհ�i̬�t-��N��)+�\���:�R}���J�0i�cR��F��䔝�����Run$�h���%�a��z�ZZ�9&j�(.�{�8.I�F/��eV��kt��Ȗ/���G.u��(�l��x��'߸��9yD� 4q�����j����d$cf*x�6��t����[��T���Z�3�8{=�?�Y�O���N�+�>�QS��0b�"?YwaD$0J�WOmC���gl3fWT����*l��#���@	G�yLО���'��t4��y��[��V@Gw�M���:e�y1rf:�����̺G�ٖ�ʨ	���&1���/�v'n��o��S�1�+�3�Ug�j��69����@��<i`ʠζT�XW�r����!R]���\��b5��wLP��u�H�	Y,f�vz�S�c\3>Y���dҴ�J��P�N�:��$�&�@9 �Ca�ҏNg�U;���ﱽ��QR�n"iŋ�C�\M.�so8���Ϻ:L��G�J�����?�����cg������u���8>T$^�"�{,�o��x��>��V��=��"a"��A&�`�I# V���:�_u��s���l�q����p�����Lcw��/��ָ��V�{�\|��c��ɢ�U�����s���i��xw���x�>���{|"�T��b��|lb͞��<�v�\ŌV�<�c�*�nd�0z�
�[���Ϧ�X�ǁ=�=��l��Վn;�=��5,���tN^�br�O� ���Sq�U�G�ӊ�lO_�&1�B�5���Sm諑��J)+��� �0d�E���8>�����)̏�yÙ8��C`�5�E�+`��70M��^����7���c�q��ސcc����w���x��Y��L�ĸ! pMn$�g��,.a;*�8Da�5�&�\�c�#��hl�dV���&�>��2և�XO�Ѷ� �X F8������/��Uc �_��x���-���LiH�����у���a��՚-�F�zj�����2�b^�0�w��D���;/".�X�4f·����"�t�1�6���+0m���_�\�����c����X���\q�H��i�ɘ$u��V@M�Lў6���+-ɩ!����8�(T��h�����$�)��4ߍ��æĺ��~�<sEQ*bzoI�q~d�nL�V2Ĳr�K{N���L�k�I�rK�9^B@A`�U&��Ok��!�N٦��o4T��_�Xt%]1��%٫������j'a�0��(9��\�2���ݳ�Y�l_Q�����h��)�
J�Sև*���O�RۛϢt��q?�ץ���e55��,�w.2Ȓ�K�i�!��_�dh	��U=G�l H��d:+�zX{߂��^�%A�*��g�������/�jZ����\Z����#0i����x'iǯc�(ܒq�<�[���و��5�:
�U����5�1"*����.=u���̪�(��_ɘ$O=u���o�=�#1�7SwD:���r]vV���+��@q���s%S�,�ɲ12E��Z�?V� ,�h�mޕ�Kø������c �k��b#,^cim�k�dpg���,�yP�������y�ŪuJ7�H�|� +H���;y�z���XqA�L��� �����֜���V+�i��f'(@;TŰ�9�ǂ=�S*��:�|�m]C��-��kܪo�8�.���.sg�A%(���FJ�YL��Be��cTb����wbC�"��r"�WmR8�cBq���J��i8vX�Q	���-������L�?{�=���?�Ә����ʋq1w}��x�/���0&�m�	�rn�M��˳��3�<&��d��i�Yi�l� "X�Ď�Y,'t3EBH�X���?̽�]Wu-<N?��˖%W!�b��g�JB�L��SzOlz	%�@h�@ !!Z��ݒlu�~����Ƙs���(�������|�9���\s�9�<ļ���ČG���PwwR��-[o�6�B�g�����.�$0����*!Lj�e9��ke#�6�<ª4O�K�.ُ&��Y�~�|���`�*��ڿ����n�|�_����ē��,<�[��2M�n��Ç>�o�t�4�c��#0%���}��Lb�'����8�mڀU�֫���l71?7�}{�cz�a�q�WK(p��6⼿x
6�8E�������ܺg�>�
FFF��g���]Fy0�G?��x�#���'>0\�c'����p��6�C�b�ik�Va�Vؾ�5�],��hps�0� �J;�6%O �dp봌��Tg	���'��O;�r�.���Jn�]���'"01D�T@����S<�^'���=GmX�R�*�3K88��+v܂�/݁�V�����\1-qe��O��]��Bi�V�trش���Y���|��k&'05Ί)ʳD��d�ԗg�˭>f�$B��Q�^r5���_��|W����iT�y/��-Z�:��0��rʴ���M�Է�aEUs�2� �ag��oE�P:C3����e���d��,+%IbԪr�){4��k�F� nI��!����Q���/7�o.�Ȅ'�"߇�����a,m�0e��<g�eX��<��XP F7~qV���u��`���s3��cfA��&�?�����z�Q�vy�Г�0���#�rV���P	�@�g�=�#�`�-i1ôH��#{�{�D����R�4��0�SY�����H�Q�fA��g�HZ=�Q��!�'�K`��4q I)Ё�y��1	�$+F��|ƥ_�
��J��uN�ѣ� ʲ��Ȇ�����|���Ԫ���d^_s�IO�:���Q�l�~�;m/���EB��3�%3�Ÿ�i��qA�X�}�	��؁�U�l�yc������l����>���%�+�ǌ��3̚�lgd#H���}e먾��֠%߶����s`b�yE)�m"8'"ȟ{��>M���Y�ּ�qb�U��*I�uW�MmV.e���Ee�lя���Af:�]�刽u�m��N<'��Fw%bG̡����s�|�^]�9�a@���L]��$G/r����
�B��z�5x_�=a�9N���%�g#����J����;�}�9�e�!�L�EhoG߻+����Y����ƃ �0��5Y&�G-�g�E�k�A��[|����Ϗ����叅���z]���<��i��8r�g(!�"��{Vi�S/�'9�r*�Eљ����]�CJ�P�?7�6<dx�;�瑑&O%���6���3L����N-�ټP淚0PBi�����{߶�_ai G_/=U�>������E�˶�=ox�p��d���J����~�ҝ^�f86��Q�r�
��U����ʷ�$4y:(��WF�o��]��Ӟ�}NX����8�"���ǔ���[��}��_B�0���!3�3?��)%��b6O�s���%(���n���*�FP����6Ţ�jA��d����I�6��.�����������l����i�aq�^���C�!ȝS��%0ܪZ���6
�Q��r�UV��vZ��:hw(���N>���b3��zC�^��/��w��ϝq���=њ����׿��� ����glĨh�:���}��7���g���w4.����W��p,�u)ѥ�q|k7l���(���T�X�[���{17=-S���2�����{0&��r�N�M|��6�ΐsD��|��d���Dyy�_��'U!	�	��[���#��t
�2::���&19:��7��,5[h�zh�g���'�4�j5�����Ip�E�f5��L�N8f���8}{Y�g;����j|�_.�l��Lk0d��k��ӎǳ��p�WcըyWI�Ƴ�\RO����߀���Oqh����������,��-U�k�^�5#8~�Z�v�����X?5)`:>V���rŐ0YX�`n��&��c�1�.�uɕ�����:�z\�_���Ok�*��/:${�$�(/d�^O��=�gdi����H=(��1A]����-���n<�����K���	�U�a��)T�����?�A��G��zV����A�ۣͦ��̠�A�>�В+٬���kW�'-9�j8@ɐ�]�U(K�^[�Q)��]���F8�il�%�k9�=������?�꿪!�H�T��N�c���2�z�t�����@�Cɬ2Pc���˛z��ʜ�5�*W�~�Hd�7����1��{��_����$�@���8�k�U;#੒��T"���~��\�����=Q,G߭�cL�ر�ij&��޴�*�M��탟_N]���8\f㹧��?��\*j��-�g��/���1Vǁ[T5��=]n4��>��d#��}h$���-qQQ��5%�\ס^��L��P`VѲ�7��ƚI���l�Hkϳ� ���؉j���+o���'�jF�dUp�y��$���,8�1���x}�z�\�k
o|����Ix��If4�N���;��~�p���<����,���+���/�}�b�$7����2��ex�k�i�Y\��&�Lo�h3Ձ�JY5,=/�'3�K���{�wp�#���
L-v����ûR�X�g��wR�أ�\E:b����$b��[K�+IQ0yg(l�F�6��"�̰��S�D@vT�0{�VOb�-)7���72rQ�U�8�Mk��e#h)ۿq�m��d    IDATeP�g��EB:�Vw�-z��)�g�8+ZO�=f�����d�=�,%i������b韠�&����Z��ҡ��k�{�REq����2��k�nݨ��<��QJ5��6{U��W%(��AM�ZV�2e�T�II���� Nh���h3���{�������ꩭ��33�����4�F��>.F���j{�۶|�3����L���kwM��~��Y��b�|e�K�9�){�`hrI�a��4��
Jq0G4����@c������-�R3�W�5��WlS3>�>T"o7[����ߢ�"G)K��CR+�_�cP #�P����W3���	+8ښ4@��ɶY��Cn(��v-�u�{����XW����_��W�\ZR�7�z�<�8�ɏ�茥>��w����7���_v֎�����;n�Ż?�U�y	��~��,�c�>�T�����xo
+�s�vK`�R��qlظ�׬V����q�;0�0Y]Ɵ�� ���c�����ڷ�nڵ�~q�r������T����&>��W�I�:L�h���nZ��}���uh��~] �Z�bj|#��,4#b���F���5�B4f���44��5}������(�p��|��W����jv
�ſ܏�����??@�V(����+�9O~8�~�v������X����M\�l��;��o��%��$L�@�$p��&0l��W�8f��;z-N�v,�r�l�Z��3bR���$�-�2������ϿzT`:=`v���fW��&��Q���?�~��k0=�A�TSŔ�F:L-b��G�k�>VNM�N$"Q�ە���U��)�:CT| u�g��rS���d*u S�[�X�T��u(��~M29{���=ͥ[b�&8��{*�FҵY
KV_X��M��{��&�K�=�K}^�+qu�����t1�y�W-�$2� i�g/#y�,�2y ��-ID3 �_kr�\�dqY�����#!$jvn[�1����R��>L��l��Wsu?c�]IƔ��[EIUϸָ�^pR�KY�d-�d�h"q��gr���!H?Kγ)����<�>f�&b 2�R�<{2�1HDO���x�e�~V�l��%�o�d���9gj-)�Ϊ7a�X�������dP&*��j_˞��G�ս��$Y��qJ�5�B��]�Xdg���O�3�Ɛn{�0����rB(r��)��-�\�~��~��d�-o��9MH��^�2��=t7��DG���!d�1�T׵b?1{� �͚T5숞�TY��i�x�l�AVޘ)*���Ͷ�s��ܖ3�����j�&�i�+�	7���y�W3���� �+����&b��=� s�_�pñpouC/��z�È3oI�G���Q��K6�GD#nG�}�k�;�����9��y'7컙�9�
����n�����+�2�4�c��y�fT��v�Jp�"�Y֒m�Q�	��Z�o{�}�n��$	�;�*���^���s�g��^D��r2�Ͼ��w���6 sNrY�)Dl��e��l�=nq�F�T�iV;BΜA����9`J�]��HDg���Z�LJ�u�*4>��9=G�|w�>a?>t���c�*sz���;����$�-��6��z�.��(��gۑ�|��\�jh�X:�G%^;A)1����'`��w S���͖��#VM��:�1m�ڙ��o��_�tl`���ߗ���Û,�#_�~u�A,��}�_�4�`f���f�#kh��V9��" �}��(܍	���*\GS�dg�#��҃g_N��N���RC�m�:���A�����Jc��J����Z)�3�J�k̄���~Q�V�D�D��y0��M�Lj�E��P��=��<����Ǻ:p������w��#Uy�C��������1�z5f��w~�K\�����!��ބ{��Y��R��ܾ��~�k��-KX�A�H&z.�Q`�{*�hJh�Xpc�0�0��O��԰e�V�y�ν�`��;$�+��Eg? /}�Y�������_��c�e�2J�5���o9*7Yʗ���_�����C�����(���*~q������;�h&З�Z	��
*J{cx�M�l6��FH�\�
����`Ŵ����j��6����f�6\�	G�������8����+��5��憨������9ha��
^�����܂	�}g����[+j �*­a	?�f	���q۝��F�i@�!����(�k�}����!�Z=�-&q�[����8z����qɉ՟�u�l��ۡ��}=@�����s�_:3��EU������O��?�9.�Ս�]�cX�cH�/å��Q)H�Fᚭ�'V��r]�T��H�iK}���9�� lƸ�J;,:�mmIoN���T˒��rDͰJ�L	=�ޓ ���F���E�}6��?.q�.iO_O��S<g\�.G"e	1��J;OX;@�Tׁs�8p�rDd[n~�ƾۚ���]��Q��]c̓Ls%�}(�(쬢k�z ���D�Ơh �U���w�6��zUܤ$�P0���D�ׅ�?�R!U����\Ƭ1!V������v��H|lݹ��4?N��U����_3#O��Y�=��������4�����ɴ�R��
��s��0sI��&0U��!�,��	�w��:�Q�Z1N�ohTR���\ްI�Ǿ�H�5�'��DR�u�X��H�;�� z�b}H�2v�d�ٚΪY���#A���nK[E\X�M�!�������Ot&��$S�8Xp����֬��i�.f1v����kĽ�)��GO���~a@:�U�:��맕ɽJ�g����A�8s�t�� ��3)�'(�j��77������ʯ�C�����#�
���WW�9�{T)x��_5^��9&[�w���eh�۪c�fLǯ��֟��Gg�ۋ�?�U�J��2��s"�>�eI����a�]�v���W��5�H�]���yj@7��je;�������������\�]��ڜ$ݢme/bJ%�v{��ݗ�zV!�WK�U��Y�o�6�ڌ	U�q�O�0?��c���ۮ�����#�vff?gX<�,3~g�9�/,��G{W䊷v�����"�پ��F�����b��k"�����D�@ǖɡ #i��>	C���5��jS)�����=�HU����g����zmb�M���|�2��J-{FV8HR���{�T��',�ِF����i�y�f���������`�w�������kwa�[B�4"9cL� lrZ��ؗe'#�CY �ڋ'.�UE��=�7"�����d!�'H����H�-�X�n����Z�Ǡ�H%`.*�J	n���(*��y@�nI�`�VF�Z��W��9�������M��xt	��"T�5�����=��=�4����buh.�q�{?�/|��y�&W���g?/���crj����[�◾���<���w������ͪ�U;���O�.b�k�:�^��N3̼�ku��@B�����%
E5C�{��8��cP�T�w�~�v�-赖0VZ�K�y0�}�Y2n�+��,��o���g�q5j�#����h6������j�i��M/�?�8Iy	?�%\~������;Z�W��:�z�(�]�:�����}�p��J�&r�\1G���ؠ��I���uϧ����A��8is����q���t<�P�O�:�W��3�X\C�λ�&6���O�c<��'`��/�񛫯í�����z�Sq���-Ӡ��� |�k�q�~�K�&q�~,:��T�M�-`��(6�ŉ�n��O9	�׭��hkV���w)z+�� �H��o��n�C3�X��P���B;�\����3\u�.,4r[��U S;��j���햼;-p���{�q%������0�`uSl5��j�/��x��b�ܔi�ؕ Ti�͞�2���UON��ԥ�I�#�(���*���D���Y��XN}�Å0�W�a� ��$���Y��X��)�'ג�����Y�s�LrH������Π 6v�C�����߈;��Y����x����U�� )\^un���M}T����-���Ex
�ä�R$�ifi��O 	#k�1&|�\'��s\�ӓ��,x�b	U`�/�y��@�bH,8	��Fr�jr#(o���=g&�p����m�$�"UG��XIG~�h
���tͿL����c���fI'�����j~�U�����X{��a��FL�EY�83�0�RӬr�J�B��}�Hz��!�u	�Z��7�� �����3� �EC~�P��.��3��+�n��u�L6��s��<t�!Ҿq0�}`Ry���v"�k�W��f3��]U@�1Y�4���Q8��y���{T����'́�UC#���F��� ���ɕ2�n���cLN&X'�Pc���ȱ9�s��;W:��Mq�sO�9v���G��<�v�i��+>2�l�k��Z�z�֦]�U��S����W���O����������=�Ѧq�o����a��!�%`���ֈ�g�5�ZC�2o��r#r4�^1�Ca��__�*���m<M�p��S�ޅ��7�Iq��\� �.!�sK;=)B<Ƭ0a��,s���10�M'�y��>Y�5�k���� =L��F6���
�c�+e5ӽ0Hл�4�z/�*�/�V,�Ƴ�-�����Zh7����v�T�j��Ѩϔ@ѽ\����(O)�X����9�NA�+a��(`�Xn�����I����L���z}��mTM����o�{^�$�.��J�'�-[7����ޥ>�����n�Ⰶ6�hs�Yp�ߙT�-����她�̱Y�~�y���==3[�x�m������=:�.��i`�xw9vN�~<�MMʔ���ay����6�;����ع�0:2^��8��X��#���9�Km.=u����d�&�1ٚ���*��Y�0M�����<К��>�4�������1䈍_�~-Vx�-l�v<���s����(������?�-\��ob�^�g?�6�y����E|�����O����$���o����I��^�J �  �[n4ln��jT�e�fl�r4�&Wa����\��xi�=�,��9g���A�\��׼�p�0�� cm��AKr"n6Qf�p0�MS������׽T����_����
�ߵ�na]��5���3Y��A����Yҕt�"����
�"��t=019��Q���܇�{L�?����|�u+!� ՗��}w���Z�[㰃��e���Spұ�p�M��ʫ~���9����d��e��q�Va�@	�����ѯ���s��LE�PR�d�ɦ�J�-`ʊ麉*�LTp��kq�=O�q�6`�^ź��1R�$�o�4���]�x�����B�.G�����0�߲_������/�Ϲ�$����$(�u�o�J����6��g��^�dO��l�"��=��i3O+��*,�7Z,�T9�C���z,*0P�pI�Ys�����&I��1�Q9�=e [`2��K��=�Q���;ƉdN��B�l~�5#0�J�m#��iNI�D?:�0� �Ep7��S$4rI�3�|�=��+���'�:h�H��{Fi�/��,F�U���ߢm/>S�"d?���I��:�����I㌨�]�3�Q��s(^nӌL�r��3���H�~��Md85P���P���	�'�W0}V�%�Fϐ��*
��%u��K`�]�4	$Pt`o��<ˢg(��=�Z���*�^1��n�.��N8�r#d��2�&�q��9���G�z�ئ��{���uVn#�W����	--S����U��� L����2��A@��ɸ*��F�>���D�tO� ��pŁ�/�V�������F����3A6���꩛YY��Wu�v��p�ֺe�=5�?���H3�C��R�d�f���6��K{��Wk�=�iV���rl�(��$^dMf�:NZo�Q/I�=�f��i��>~�.�����X _�m�/)xE��H}I�����@u�:���i��z)��$Y�6�z�T����YhV��Z�2�-_v�^��V�7��1��0�5�{��J �c����^J���;vY��"TIg�@9[q؉��}��1k��4:Uh�eߒ\�Aب��}�Av(;����sA�;B�a�hk�`[�a���`|-D\��sx@�����Al���&� tHR	0���VM�S*���#{��]� �H��@��Ggy����P�P�ls�����6�\ʽ�}_�VN�-�jUI���W��e��+�O�Tj���e, F�vCg��$�����gl��X�b7W*�E|]�����p�g���~��n�|��n�.wİ����D�7�r�R^�1�i,OF��hZN�>�-�c���͜�?t�Z�9�U�r�)x����^�B����Q���~����'���vBudTr�-���>�oǶ�'�_(㚛v�G��sK=���Ȩ٣��j��7F�υ)27'G��1?3�A��~�}q�럃���U��l����VM`�j��4�y��~_��7�o��+��^<�>ǉ� �y��ǿ��]{�\y�%QR�v��j43�fN��Z���)+��?8R�a��ذ~5�&&q������X@���>
/xƙZ04/��Ux�[?�����(W��S��kh6���0�Nc��FK���>�;�1�����&���p��&��q>Q�Q1��]ULi��US.���(�WM
�6�tk)�R�M�$�;����F�3��6U��O��;�z\%\~�!��_��C]s$��LJ��.cr��vcӇ��T)`b��S#x���'>����$՗�kص�a���@M�v@p�8l�\h�Rl��t�X�&*8f����w�	����H�׭��a��d8�tzvK��E�*����6|���q��9�~���kVLSz�>',�1y���_՜��7�(v38X���@���c�nh8#ʀZe`%A������8~�$��3�$��5 ӡ@E%��� A����σ�$������� [o���Fv�X.féyM1р�J���F|�2>�1O��&3J��}#yO���n����P���p.p�4ɒ2�C��I����d�e�h��
�ل>��t��I�{�,aw9d��c��Y`T�����"Ǯ��%'[�m�qST���UO&�\F}['�9�=��#��{g�y��} �/�V,�
D�0�u��U�l���E�M�T�k�tv0�7b=�,N����� &]�Bi�]��Ӯl��J���HpN>~�Jb����,�]�U�j��('�������������]��O�ɥ}K�W�=>7�w���_F�n��¼(�ǂn���%�AfEL�K)m� ���15�[�a���g$U�|c��WT���ںI�&^?U�'9��,�0�q��Ƹ��t^�b���^3���죂���pC"����l�X����817���"D�W����z�g��g\�z3b'�g�X�xb��9��?�؜B���2(��o�������ʼ��=��~��ї�,�lf����y&��z�u���ʑ�AT�.H&q9���zL��x?�L��ͷ�3y+ל47��D9q���D��J���bRAL���z�?��}�����ۈ�T��=�9��,��Ʌ؈� �S$�����j��3�~�,�y!�o�n�8���,F�rt%	�4�-a;�GA
�2�(���F�eɔ�PA��Wa�RYJ�� �4O>#a(��mw�g��I�ej�`䙿Y���s'��\<�i߹�S S:0ma�;��?�4��/�5�����p8�SR����kwc~PCkX1M��sM�*���1���*5,��UF��v���Vo7?��N{a��j�S�Ǜ=$(]�9Rcf?�O /z�c��= ��m�%OJ�/���%��o_�f���Y��=�18���zm������ß�&v�_B�R��g_*)�r�0gc��?��7��X��Eo� �����L�#0������t6���|�&|����e?�FJ|��½�Hc�    IDAT�Y����m����_�8�ƀ�@�Q�n0� dK�R:�4b��$�,� &�m.Y�P�U�i�zLN�`�Z��=q�7I�;R��k_�X<��B�hr��X�k��I:L�
g���j�*����j�\^���T��b�0^������?#L�������Yܼ��6Fe|S�U�Li(3h����ç��X��>6���qm�F��Rm�Et�S��b��~S�gL?��w��&<�(�;���o�4��cdlB,N�ʑ7@��@���^��~o���7��Qg�����ؼ����l�����߸���eJ�9��Pm� �y8ꈠ��J���rׁi�Fq��O���b��(6m\�y���g5�����[��fg�C��hv�h�Yh�q˝".����gW��ᆀ)+��$�5�ġ茦6
��\��3�*	�ce.�ݪrJe��E00���͓��d�H��������6���5�:)E��0x�6�e�4E�V#��J��{�J��� |qRB?`e��Xga$,��KB����؀B<��Qr��qf��)�����~�À ����69�S�-9+�*��$��dؒ*�_��㇮�¶Bň��z�R �\��A	�BW������jr�#����P����uJ�RE#2Si��}����V��N��x�J�ӆ��\b�����+Yu�+���ߑ���$.[�sŻ-�U��ד����2�0%|a$�����ӞG$�V�0��n�����|�v������V����s��;;���]���WL��L��EC�+>3�\偩_�J���O��
���AZ��Ք��{�Z$����f~f�I���x�l^��#�Q����d0d�1���HQ����k�Is&�lLf�9�1�C�*H���7��k	�F7�B��F&�Y�h�i�C��ճ����+1�Ȯ�����V��D�p̌*�Td�S�S�7�|yWf���O�['�ݤ��Z��l��q�}�s_v]�ejIy=F�k�
/�/���CsqO�4⣏�҇��㤕E��48�є9��}���z�=�D��*��\�b(T��I!�3��٩��x��D֝(#�əJ	�!�km�f_�%�A���򼌹����}4aDxX�|����<w����m'����6����b���|��^/%�����>K�y�__��?ڼ @忿��1��7+�T��}��38��3Pٶ�ʛ6�\�#7M�(�b���l}�U��ZJ�#kO�/�q�PTdkH���tk���О�$;����S�6��&���8������a���s�}
���p�\�軸�}��W�F6#�R�`k���;�J�Ky��c�?O��Ds�Uk|N�	+|9�3�}1����d)���sL8;��e]o���Q�?u�����9�
b�Y�ݹ����Zܾs7p�ix胶c�l�k�_ݴ�����MP,�1>9�5s�E�L<IfŏK��U�v���-��3�����>k�����"��m���P~��.�����ҟ]���v��o��?��l(b��u�[8�#_��7̠Y��U�Z^��bj7�$���*�5�Ԃ��<����I��}��;w��<���Ɨ=�;�A������x��}
3<��P.�111�Y���X�Es�JX@�{/x�c��s��x����nk���4n��ٗc�sCp\M��]��TyW3����nVL9ô�jc��@�O`mO^�������؋Ro[֗���_��N�нS���;�Wo�8��Q_%�%7��{M�ֆ�����/}ޓq��ը�A+v�o�߽�Z��\�=�)e�)�x��fR�ð�Fq�E��A���ԈUL�FK�v�Q8m�	8j��޴k��MF��"(�X=Y��l���[&��߭��czf	���=2|Ut^���\�_�	T˲�ʱEl�0�~�`�s���C�F��%A�O2�6�MN��D��(�!�����e���^�y�J�I�ĀEIJ��>:[BG��93;8�)ҠB���1��3�Y�E*�}w����l>ɟ|e��Zj����\�"���1wY1���J��(U��R������!M��jb�)-!���rY���3ƚ��I�lZ��� ��g�*�������#�i$��7u�dՎ�����0����z^^���9θ~8�8�b�!���'N>�|�.�&�gI)/Sr�\Bf$GQIL&=4��2�d�/�d^Ʀ{(%F�.E�z2�{蚪�68�n�6�pxbf��]dS�4���Ki����;)_���3\02�H��F�������XTM��
`bqɥ�z:ߺ{f��;�����	�Ͼ���͸a��\��\à&�
�Yrt���m_x���%�wq�G�J��L&�;k#��v�o���,����yˏ�3�,�f'���jk�}.�=��/̜"U��X=K��0˪\C�fRK�+s=�(V�}�
Z���U�k��#��#>�a0��؜����i�n�k�nl,�G�P�'Ʃ�~��d@�M��E��ALY�k,2��6�ˁfD��M��)i��<S%�3`ủ�(��IlnVn�hm�����ŗx��YCK���ͮO�lS;Rk�/z������ɛ�[2��E�s$������0y��WjY�J�eJ� 	��e1 SX0.Ƕ�T�� �D2����v�K�<m��-D=��!�3trR#�)��)Pc�'�_�K���:ˍ�p�yd�*��<c�1Sr����@t�	���Y�ql����QI��*�S�0���޶@�1�͐��:0�tZ�[����@���G����]��>{Lo?��.�O���Ø�V��ntg���#�0�|KDQ������� <(5��сARcQ����g/�5��X�G���A�0�3��_��y��P��ʷ=xh�NW�kl��MM��9`�w���im��7Pۗ��w]�7@�4���	T�FPఠX�t@�5U�"0�v�47���A<����^�tL�4�3�UB��O��l���h��_q��i7�����o~��~��9���ٖ��[����97��G�6�8sA1Z��r.��#���f�S.���2�����}�V�3x�yO�s�~�6E{|�[��o�,w�(��Q*�Y9��K`Z406�A�?���p���gaM� 	�U�zx�?�kw.�W�Pujd|��&1R��̝�`��D6�R�rE�����ڴ��9�JE#j��e,����}���e}~�=�ۉ��wt��Ww�/_�!�`d��҆�suj �r��գC<��w��y,N߾�����9���#\|��Xl��+��?(�T�#�����r��*�m�^��[A�G�X3V�h���7��]Oڊm���7�ú5�Pg��w��\	����F��+�*!�dw~������x;�2�:C4�Eܱ������]�P��j)��o�4�t�fA^N��Z|�GU�x`iiQ3�؋A��?&zV%bJi<`s�tHh�"���l)���:�aa�)(�cX���&I�g�Df�?L���0�1)���n�a�*�]2�� �:� ;x	#�#�c.-Y1 =��=���	
-��2�2�fZ	Tfj�D"T�ٙ3`�f}b
٦����֏�<���k�R��O���I�en�	N�f-�!)����$|�br�t�� ���"ϊgd_��H�!�w���x��=��:i�U#�a�p��0cOzS"�Iǲu��_���pF50K��F��=r)�̭�#�NG���Z��=��E��E�N�X�O�W?GCJ����3����Z��[g.�My���Q5�$�����k=�S��Q��/.Y��k�%�UU��J}|B%�����F�[�f�u�UH����q4�N=���tc-�07��+nH�Cf�{ӪxaX�Rz*���v���C�{�w*�q��R�UY\y��I,����S�g�>ŭH�s}�u�7����,�N��窭+�
��v_�a��/���	]�#��k悛�oM�[���ci�P	r'ɧW�IU#^䈣D
��������]�)�o��A	`1��֒#��x����l|DF��9q�����r� �	���[��@"*��&�}�)t��˕\aQ�L�=�θ���{�{��7�o�H��z��c�&^!ֿ�_��7H"�1��w��T5US���`ha�G�{]9Lр���v�YZF���t^s���5c#�T���8@�J�ˊ;�D�RZP�PU�ӱi&l)q����Y�y{�f
hfJ>�I{� �������+[�سZ4Qo�K��#���{��T�X�Z_yT���7����m��9���	���Rf�L�Mcm��:c�mB����nH 0����0[|�ue�h���<?���<�i���)����ၧ�WC0�t���?{~s��x�#�£y&��(ٝ�o`�V��xE��%,�q�2�束ǎ��T���jT&F�>X��K(��ܔAeoN����r{/y��q��qsP�Rػ�֭�x�ή�`��CC��u��5�����;q�1S���?���T/�3w���O���.,�G0��!��j���`�M�������C:6:* ǅ\���` il��Bc��%�< �Zӷ���8�	���.������o?�V���ZF�R���4?t�P+/c����>�,���g`�Ω��5{�ל�	\�s����*&VM⨣6ar|\=�2`�d�U8>Υ�2����( �f�aV�KoC)����(�g�yp�'ߋ{�e��2��_���ؽoc�k�Y,��@��j���ZO��/x��p�S6b���{��}?���iV��.�XS�p�h�Z	��[�X���ðז�RaH�.&jLV��b[7L	��r��p����a�Fh����]Ҵ�Q���oo�����̅�[2���ob�a�K��"�=�,�p��w��?��O/�7��u}������{�XW& ��)��Y��P���I��q�#�J��oJ�?�|�Ʋ:�>s�&����
*��nVN[UNi��EF]�x�5��$)�88}d��9Ó,�f2*�^IRP�d�e0n�p��%��!'sKF�*����p����'v�X �8h�BN��V�l}U��5}^��0����Y�+�A���<{k�H�8�~3?㣤j��dHڃuNy�'�fӒ�
����fGI����&�c�b?���IϏ�!˪.Y�cM,Qv����rdO�}k+�����}e)���͐Kr%�ˈ`%��dP�ٌ�����)��U�3*e��J��t��7-Qw�'����m��x�beq�� ��~Q��v֋l��PM�,�xL
�kP�(�X�y�[�\'��6ʿ&IϪ*�o�e���ϐV�sZ���I���KV]p�H��ST��U1��0�����k��JF�YL�����J����r��O`�dۑϺ4?��m� �u}�Y��W)B��E����b��QI��d�;#\�zrն
D�Y�^���i�`�b��ڳ���11qW�;�9S�x���9'`��w�Z�9��s��NJ+i����F��1(�<�$��1+����>��r��K�Rp6�ʝ��5R�G���4�_v�����߉���*��-c[H	������ɨ�����}���s�ܾ���[�#�!��h�'���I�<b���,��������K]��zӝ<c�{��0��Y�թ�� �
�)����B��Ro�A��~��vcY�D:#JE��5�jUMP�ԌoT�	叽O�2:��Ub�#�8�2g���x�%5��C_9uق��R��s���8ŔӢ�X�nG�t�7��:�1x�cNńSM=ȭ��f)���Ƈ.���cK�t�UI/MB�)�V��
�g*)�7�;0�O���2�UJ�-U�vʜ~c�ۼÐ����٥|�����,�a�<�����~��qߓ�H���w��<�y����o�Ӟ���o^���G���	z���Ƕ��������-������������5)���́у��vS��a��ڝ�߼�qx�NGݥ��q���~��N<����b���Zx��x�{��˯��3����y��E�x�����������R�0LY�`�xx���b�����[(͆�Iz}�Ґ--��ca�0
�6
�x�yO�3�thV���x�[>��6��ɜhdtޟRQ��U�U%�Wx�9����)��� �xx��įo��R��B��ѱ	lذ�׬�X}uV�|�3<4��>�C�����0VV2�
j�jl�ѕw��i����c|�3�=N\e�^������_����Ī5k�j�:�]��s �\�k���pϻn�S��8��I�����补���W��/�wNwqx��~a�bh+5T�2+�v4h���L���A�@�k#�&k��kǱ���qʶ�8���z�&L�T����H.䇎��8~����﷿�aVA���q����R�.A{��!�}�=�����Z��V4:D�4D#���L.]�H��S��9~��-�߈�'^�"��ީ����l�7���͠�/%2�$dܜ��PIڐ���z�)�-v��G�4����dRĊ5��#r֐��J�ŕ�H?��-i�d�ek�¦���bƒ�yF^���*�&�	p��
��7f���*���5�Lx˭�HtHd��JF�SI�Hj�r��R��\@�3x�����@#���U�t��Y��h�Q��Ĩ����cU�\�ճ���O��ɛ%��e�9!���l�lʁ�ea��+I#N��Z�e�f��[XV����kf"aP�%���7�?�9�=KR3R7����&�>C$�b�ErX����&��fi1�G���h���o��f0|59���j3eU�p�֗�Yd��ٳ������A�{� s�����L�Z��]GܝH���?��7W��59�2��׍?m=�ȕ�}�	w8�T�s�<xWC`jk&�f=6�,9`�5~6Ε��E���>���&�G-MT"�˪'��,���t��u���=��M9�ⱃݘ��Ki�B����Gϱ�b���֑��0EPr�"%��uX[@�dH/�� �E���Ϙf���Y���ې�+Nj�T��R'3�R�>'�W1�?�I)��`����<��}�=�w���ҹ�UW����o$(���F��5x5�kQ�'�|�|���l�@Tvs�[�aV�t��OF~ٟ�5���=���R){����F�)<��fnL��+�//��*���@�g�b�7:�IW�^Xz�D�k������(x�L	jN����̈�$�Y)mqjE[���V�6�7J�"I{SUFH�AH�?��@�3�r#���b�-	/Պu�:�\�c�&�W���S���0�"P�����V���nm���U�~,�yֶ��bi�t���W�v���p͝�X��!0��b%�$G:��8FF�ŷza�r��8�����$ْ��?�ߝ�J�=0����OFs~��8��x�[�ý��Rō��W_{���`��x�#������~�zU�(�|�?���E���/æ5������w�����	W\���8�V�1�������Uy��JSo�B�^��Bs�{��xң��^������+�F��ƽNۆ׽��ضu\}�O_��-���/���x��g<�t�j����p�u3x�/��C�`�U$nxVn��#0��eTK4���U=�!�6O�~n�V��9��]���xՋ���@�1�Ӹ�Y|�������'P��,�(`z~	��<���^u��ǟ���$�`x�������K4���UP��att����\�Z�̤�Xl5pxn��K�̶���j�*<��-�w'f�A����H����cFu�5#���7�Y�%�7�X�Mߺ�gX�f5μ�)�8	�s�� ��u��Y�m W�z ���u��7any�Be��R�R3@`�7���sVNKE>�.��&��6�+����Mk���͸�	�`��[�a??a?�|����;����9\i���(+ow���D�C�*�}�4��oq�-{��_\���g�/�0���:uzŅ�I��fq`���ꏝ��,�ƞ`U=1*B�    IDAT��֑��5��/�9��ZY��BL��܇ok���=˥A�A�VG���m0�3�*IҌ�GG��h�^�}{��b2�O��~��Ҟ�'��0����j?iɵ}?U�T�'�Hs��=R��g�%&:?�-�V~��H�L}k�] ]�e$�a�dy�$|��X1�{o�D3��j�z"��Qxe+U��(�H%���Oq"6�po�{R�"�
e�H6��خ?K0�
��`[^F�����i��� 9s�Ԁvk<T�z��7��
�@�'��$ �V�K�s��,�u��˲=�MUi/�/n�qE���ШD�*+�hcĆkg������7��a+�bV9RA=�Ԣ��9C6�!���B]
�ɒ-���i8S��l1����"I�c[zu:=^��IJ3vȣBT��w{8�[V�w�ߡJ�J�+#}���T�s�.Ϯ5S:���&eY�3f�t���z𒤝�rs��,[+3�gJA�y�1�B������=w�\����P2�2#0_XUsGf��9� P��/"���=�:@�b����q��z��ȗ�<�?C��&�5�3U������� ��|�8��Z'���c�БUO��z���Y�bX�������7cc��;�J�*>�yN�\s����sj[�qrF�6e ш�\�j~��NO/�Ȩ���R()tV����r=��Q�~Z��d
HW~A�Rv��3t��S���>��cd�
2��#kE�|��h�}W�+����q� ����R�j��S��<��E)&�Oy�8����۶���)[6��12=�����e���I0s�\�\yMr�+����+v1ٛ�k^�d<��[A�%s�#�=�[�}����_�]�P�J#��j�u@� VK�싱!�v�ù�:�*uN�ܐ9��/�@RT|a���n�ֵ��VL�s�,�}N݄����ǉzVD��f<��/���{�г����oqʉ���|���&������ �N�ލ��x��?�_^���8Ƨֹn�����>c8��z8Ǵۢ��@v�ݥCx��'>�L�\s����{/��i��r�S��?
w=q���-{������8牏���A�.zLy}�f�7��"\s���:���5����t}��P�u&�Q��k���M���m�P�����z8�����1m��u%��{������C]���?�����y-^�����6h��+�W�l�u��v�r��te��uUh��5# �E�{=4��t�3 ��\��0-v;X�9��z�/aU��?�>����e���G�U�bQn���ZԺ��S��1��br�4�cy\v}���[�y�,�}�YZ����^�[Y+y�
=�t#�V���45�c6���'�{��[�Z���:�5c���������{`�������DI�r�+ �^s�f��>0�_\y#��y7�I����qo@#��o�HU4el�׹tE��A,����\iJ���nV�d��$���g\�h����`U��)��!�+S�#�?cN�m=�d�%#��l�ZV?+G��z]Y��ܙP7��֙�`��s�7�oFR�H���[Ƀ'�|F��z�����eY�.3��d��&8�9-Z�T>9�����\&��l3��P�ʢ����)E��%��p��f��\��.3;�_V8\ZŘ	N������Ğ�i�@L�����LS�HIOT���_H��6��Rߍ�����N�(�Sr9h$�l����FT�d��4�=��@{'��V�����E�).��V�>����MB�ՋX������N�x��f 9�� �1�2d�+��5U�-��-��p�!�j��G���M@�>O�YE�x%�)��1~�"�K��������G�3�AP��;%�9 �5m2�LJ�x��R2�,be�J6��gC��4d��|r��=�Lʽ�U���<6�,׫�$���@�?&�^{3�e���\CVQL�2B7sc�T2J�ۉ1dX�|!ک�|�f$�[sZa�o��|\Ng���ȍ�LГC�G��./�Nq&�ͧ�r`�%�;�z"F�x������mN����H������G���{����+��o�v���aJ�8�t����"��s�|��i���@�H����D�=w��13�7�ƙ8(M����X_	?�+̰BYf��{��x�GSD8.SJ��d=�$%�W��F<��x���
K���sJ�j?��FG��PUR��X��1O�+�(����.��(��R�:lGy�����7�	�� �������yfxXM)�*��
����g�O�b
�,����O��d;�o��,^��O��Y��'�Lw�v��������\E����Iyc��+%�1�O�@���M�S@�ZC�cA*V�
���m��j6]N="�d�iF~#�����OBoi���8㮛����0�Ù��e����s��^<����~�q�V��K��v>���F<���)�H=0��n>��_��S���=(U'L��.�j��n?B?�����.�E3 t�p�	lݴV�B˭��.a��F�þC�i��w;�$lٺӋ-<tXcKN۶O~��v��K@�ܸ�����q�,��:�X��R���X�c.�^�SF���JVF�&��^�A�a��%�u�����UT(��;��Hu�R�������o��s���bU(z��/����o݈�}��h�'�pt�Hט�D��3(�R��r�\����}�����;M,L�G�1��r{�[����7}�Q S�4�٥��� �q�a}�S�_����ͳ7���%����?~�޼_�^�Aj_���H�E�r�la�E�Ow�!����)��f�������'lـ��&�z��u�2p�?4��9S �� l�wsd�$B��M,..����+`�W��rӍ���6\y��wx�b�!��8F�p$mV:�̈�$�qP�6��M�����);�P�)�;��F�?9�����o��h���-�H�NO&r�e���zy��pj�S��%�p��x�-2T�َ��z�٩J�X$%�W�2������D.Ⱥ#z��C2�9�J�D{���p;�}�K0����^Q׫YU6�`璵8�����)i߬�/�3g�-F����?ok�p����T�`�s+�'�뇠�G%����k5C��K��������%�O~|I:��=y"o-�H�yv��*�����u8�+K�m���i�,
�Ч{�'��a�$@�C;��kk��c��NO0���?ß�d5b�����L���"��&:�8{�[����=�r�F������u&���G"�ĵ��$�7/��|�_���f��s�L�`;$�/����ND��?��L	f�lʋ�)���&���de1��!F��*ӝǋ֧��^i��l��A2�}�@��&ɡ�?�N�=�:��q�*�^�d��<-��c.���N�b���i�����������TM��D:T'j50 n�L��U��ǞО!yc5�Ї�X�v���"�زQ�%쩒���������G���3��;q� ƌH�����'/7w�bF�e�?T=&�%;�;*����*�s	?���� L�<��5yqT����)@��qC��@�^�����N,�<Y=���B}��؞�ؕU3��>��!�*�e�dsn��/xxL����UD�j(7�R�0�J�l.���^��RS�=Ls]6$]��������2:�8��49j��c�b���)���Fz�M8��M!S�n�)�����
7I%���xY8����`��j���<���d��yy(���9bgi��v�A����))�_�4<�~��RQŔ���)��W�r �wp����1�9��I��S��='�h����1dX��ּbj,�^��V��N�����nQdZg?�}n{t*��\�GgaVf7g�̊�y��q#��n��K~�+�{�+��!�����=���6Ҕ������v�iO~���P�Vd�sˡ^����k�
���bŴ�E{�b�� ֛�G���żpTH��-%���P���s�9����F�p�H���>`c�"NںVOb|tL�w�����p˞y��5�4�aW��=�>_�b��94���_}&�����O�?�S������Bl��H���=L�w�g�&���˰i�z<���e_!�^rm�·p�y4����"I��	BB�q1���:������%�w�sYi�Cgy��iT�x�S����C�i5�I
�pw�
��K=�����.E���#ϼ?��cU��P��g�`d`�\|�A��W��3]�����˴>8��a���5-z��;(;�z��8z�8�r�Q��	G��c7a��UX�f*5SD�*������ l��K�~�67x��M�B����R�N_r�v�!/�q��Y\����7�f�+���2�T&�6G^1�q�xB�X�D]�
j�m��q(η;k���zФ>_���\Kr�s��ɲS�1Nf�H"CFҀ)�$�
�
���f��$�8���"d�� y��1��l��AƤÁi0���z;C2Wp�U�*@������hHk��~�c� �[���l	��� �jg�-o��8��te�W+X����Z�U��҅Y9+Ȍ ��������,z��PG�"�v�R���� P��i�:��h%>G�� (9ͩMl�ƈ�~}L�8Y%�	ʽ��fD�}êO���He�e�q � رvx�7ي
������?+A� �'���'h�g��=9=��x~Q!T� � ��Z�袏.3�17O��%�12+�V���P�*��!9)���zu-�r �"���!�{���\{�v�������g�\ L���.�Z	P�c�Y�o냏���?�5�9z�����Z�9�c�����'����o�ٞ�����=��<�����Of���l�y�|����i_.)����(ֳ�Hm٤oS�f�G0,E���@���גN���r�Y=?'90S �`nq��g,�X�������\hJ�|NZ��rec�e����ѹ�4$b���{��S$Κ���8�)z6�6*_#�����֋ hFx��`/���:a�b}����3��M��5���J��9o�)N�"����{Pe���F'��(��p�-�F<>�>W�)�H����M��y]�({�W1��N����n���􈤯Ib-w���I�rQ>7f���@��^��~��Dt��>a�TuѬQ�a|R��)=4۵����M�N|��hDkc
�����	�9���
�m;��)*�2E���L����lK���B���Q���?�7�����mI���bJ`��փ��W��,c	uڷЫ-� �)���F�'���YL��Z*k�'�:�8������v �,]0 
�ta�WL�ٜ�F�5�3N9
�}�y8uk]�� �翼
/~�+�{�<������5��-*�����W��V/�Kp��'�r�1����ſ�	��F�֣X'��hEH�1e��{;Y������~��x (�P��/2�x��=�{��-]X�����%r|���q�j#(��(���T�~��i�۴޴Ὂ���l^r��=�F�eZsXUk�YO~$t��X;Q��1G��w��)߂@�2��6�s����Kp�Q���zK<���������	��0(�$E�� �Vp������l��V|M!���G{	��C���+�11R�7a�1�`�����D��=�Y��7܂��tmc�2֯���SX=9�:�����X�`���M;��}sXhqn��U46�E��frU�rʊ4�r��@�t�^F�S@�m�U�X7Y��'�{�z��XLM��R-�R)�*R�A����*Q	��o��K>����:ټV��N������D��@�a�7q띇q��p��w`�ˇ?���@)�ג��-�=�q	�$�ؼ�֪��@�~(�m��p��?i�E�P�99>H�_Y��8'SL["S�R�Nh�m�K�^��� ��#������
��YE0�3�n��؋��b�lm/d����}~�6F���3ƒ܀����.L�Y���*��%1��Ǥ��A�'�kB|������$�ai>a�$ד��8}N'�2'T{Ѩؤ
�f��)�I2�����o�%�VI�!V?�-.g�җ�q���-Y8GfxU,j$�oϞM��e +�gg>�4GTd�.]��R���Zn�{��V2�Aڹb#�Q����6���3ף�Dۚ���{����,�g�>�����%P�\��̈�>C�Gq�$zz��?��r<WE�dTr-��* �~:ˬ2�8����{�x��ǚD�+�B��;&�\����gl�6�Q#B:�{���r,GTጵȀgV%�Y�k��'F21��ϻ'�>��.4�!�2sI��bϝ��~�{��e\�Z<!����E�1�ť� *�&�eo�5X�D4ߛ9�EO~�[��	��Q6c�~�6;��!Jl�lVl"��`�b�=� ]Vy1ZĮ5���n?��X��\U��ٶR,(w�8o�E������To��;�#|FHe=��(⡞SH��-�6�^'�f�he�Ԫ�4�*�}�R���ܥ6#^㞦��$�T�RCr|ӈr���j'A���,_�SWX\�]�kE�D�`?��}���T�RV\��� "��",}|���}��]���Q��Q�>b-*��6��z1I�8�
)���|F���ƶ���(��w���oh���=��*�47"���X-eEV���[*H{D�^�%�����-���.�jE�Z��='¥W���MJ v��Ȱ���<^������Y���Pȕw�p8�ͭ�}��]D�8�n��n�����sg^k�7� wJ)?�,Ϳ�!����O&ub��ؕX$
:�3T.�q��t���87�+����.�^��7&Y��}����O}��x���g���B�"���w�7�Ë��3�a�l�z^��/�k��ʣ�0�j��� �$�NN�#U�\>tg5�x��9r�v�;���hIyo�k����3�Y4_/�4�KC�P�M��ߵ�7�(Kd��o�0�� �ugj,����iO�	t�0V�a�TG�����UY6e�Ue��(��bvq7�z;v�9��IV�ƪ�1���QR�7������ /�Q��J5U�T�J�RQU�!����O&��fvm��}��?�}ٯ�[V��k����9�ܶ�(��H��J# �AKb�&!Ѩ���"�l�X�E� bH��%h�y D,(n5ԭ��n7�_�����P�r�4{5����9����1v�Z]>����V�ߨ��Ҳu����dƲh<W �=Ro$V "aPW�Z��YĤ�3dF1/�w��ŭ����`�)�j�/��h��X� �Xofxq հ	M�����w�'��oy���s>���+������:]�Qo�L�'Ӛ�u:_p܏c��M��q9f��Z���o��nH8�Q�!�F��N8����^~�q}�o�o}��;y�^�]��tdQeY?�)@)emnB�X��T-�/���c�&P4����G�^JK�%865O���A*9fP����MB绪#d6 ���^kx5��Q�O���%zMd�	�q��SOGA��ɒ� O�N����
������
 ��u����&�o�d���Q&	�%�&駁Fj�RӘ��Z,��2y�
^Z=�7q2���Z265�-�#I2�<��%�p�˵�{I��E�4��d2f����&&�$k :�y ���;�k�i�mo�zJ�2��aێ�᧱K:=���в7�#A9����=��i�՞�R��KA��2�=T�yg�E�ד�A��qMa]g$��Gv�C��۹�t_��W�ޛ����a�� F�~x=�� <��`Mv(RyG�;�&?c���
h�h�6U��u�h+�����{��w�OH�� �2��Flt�+5�� j0~i���x�k�W˱�D2���]'-ip�b��bg�s�ذ�A�bE��    IDATE�~yr��O�W��zg N�G� �-��%������ �(�a��<�?>72[�1R��P��a�E3J%V���qD��t#��LMo�$���E ��c=�Bh�\?Wfys^B:�2��o$n��ʥ"mi�9���Ib)�$F��G�D��~ Ş��6' �SR���=VU�ZQ��#�B���ӻ�|��h`*ߠ��!�8zPM][��d^�6PT!^��>yw�'1��	곣g��4*�*^�$6�;~Α��^_���&{�]����Zf� Պ�	}/�CR�`��،�1��ITڑ�l���DB��7��������l�|���#��0MLQ�q1Oף������]_��-cJr���h����3�X��q-'g�F~'2�)�iv�W�Sl���x��6�)���l�+��b�Ę�J֡4�Q��ù,N�Y_�ţ���~T�����/x��������>��#tخ�/�Ywn�1Ӈ�	��:����_�/��ϫ/���!RW������Z���ɪ9 �s5���d:3`�35�<x���4��M�@������7T�C��Y�!E }1�R.���R\�z0��iJU�3ϡɣV�J�D�E�"�u cp�d�^m����!x�#�^bG'�)���aA�����нCL禲f��<MkrZ��3����������G >�t<�Vu�� �oȨ�; ��i����,i�(_���|^'X�g��	�-�-�X��Y/��T�P�/��Gu2_�٭;s���N�!.���"%t��;3�0 304�]M��Z�k~����n������0��.���jv���zH�P��,���Ϊp��W��-3�L{[dʴLjs@�[�
3K�G���U}�W��|�c��K����.k�G~3���u���2�U�9�q�i�l'Zz�w(�� p	He}��l��HҢ�nE�R;03e�B-�m� �.X����ě R�S�$�{fŚS(9Bd8ڐ���xx�ݎI3�}�U۵��Q��/��&ұ8�{�&��o.wn��M�0�=�"Ǖ`L%;0���R:���T��hmv{:�hD0�P���{75яM���i��Qj�`�7��Ed��J��;�7��N���u�	_�����;V)���O��5�|b&P�^�S�0��� @���!@�3��,6��d��l���t(���ď�ׯ��5���6�x�`5��K�� �#��/��y}��\��D�?c�t�������m"���reV� 6��l5b�ًMh$D���3ݐ���z4�r-�2�Vr�;��I�q�s��%�������(�Ll��Y��δ/�Ad�/�Nq�*返���h��C�iq_�d���r��@I�_���&�^2���d?�	|ɞ�{(JrN���'�Ne��9��J��+3,2-q�2�9p�Q�u캚f�wQ� ���dv���F%$p���{�d?eO���hC����~�=#i ������R�>~���#�=��j��q���GB[Cu��s�Fr�Z��~h�Q���r��d�(3ُ^@o�:��2�����X��V����9�gC~p�.���o$�%��/�NT~x!Q�a�6��#l����� ��D���0Eڳ�޵�#!����Dr�@|7k*� �e�����9s� M�'�-�:�f6Y.E ��p�f�����tn�����B��		%�y�Ӱ�R{PM�Zo�L'�C#���͏n������o���/��P�⭞�q�p峑1���R?��R��ü��c�1�PbB�G���GX2�8�)2Z[��DaQ�1��^�w�dj��)�`�P�tuz~J������\�����ϼ[�����ԗ<ۚ�`�I﷉.�����Ї?T���;S���z�@�¯߯���Q��g�h~��l�sM�g<����➏����"`�w��"p��dc+������f<� O����Y
�ZR˃*I	��e2�Y�I�m4���["��]�ѕCun�8�Vl��]/����@�v2��ՑT86P����$X���n��!B�wB��*@���2���>4���a������5���^4	pDV� �,�)k�j�A�00c�sZ~MJ��	�1t�G�u<�O���sW3���H�wq�"��av�����dW��}���|v��������g��z��O��?Swn����{*L?�ͨIm�� �N��&�T�@���^{pU{�~��>R���W��X��qdz�hh��;�(�ym�>vz�(���D��1+�%9��e+J���cܟ�]*�l����h�)d.�,� �9ãdQ��UG��)�N��:��?!.Ē�{�ܗ����&R��{�|ˌ��;
��Ƴ���2�>(t��`�و��@�Sn��w�n�d��~*%����b��ېE��NVɵ[�(���j��������]��dA� ��R�6V �C�4o�G�7��o@&]��)`s0:��-��Or&�@�nã_g���T=;��0�&��=�@���˰�d��.v�AVC�4�	vξ	�z�����~���K��rI���q47dɳ��N�`Q�t���}�] �7�SY�c�gǸ"���up�+	�#>̱�>�)6�
+��Q��a������I���H�w�Z��>�\o�����c�[� m��8%�#���&K���=������n� �Is���\��	"jR�j勳���<���]#mߜ�� ��]i n���UL`��X����Z���!��u儮YM���W���GdOzs$��8������!'�h@\���X�������8�P���%�W3��ᨠRF��Q��ߏ	��T���ڈ �Rsl��.���D�񜉽��$Sm�ߗ?�b�,E���ㄢ�=C"��DQ�M;QT$Ci�X&T��q+Gu�C��͘:�jMS#���Zp�O�>�FB����S����tƩ�� ��͒��!~_� ������ѓ	)�l�Uq�����)%9�u���fG�_�Q{5����v��M��n���d����x�
�
q6@)2���U�._��__?�]�R^4�CkLL�ŗ�����w_����ZAʪ^���L�9��!��R�h��Ҍ�'F�-mҵ���!�A��,����(:ͱfK����)k1���z����Z�x~Q���r��o��^%>��p�ѯ�U����������x��������_���ڎ�9�����?��ڟܩ��Nm���b^%��E�t9�3��5���95_�O�cx[C�R��!� HS�&�3�'px`����&��yl ��a���L)�����u2ؖ�jSI����e�"x~���
�s�{}!%�f@c�x�|M�yF�%�)Ѡ;� �|cbihD��5��L0mPp�+�S͛ &2�|�G0Y�7�� ���z~�^�'�qaĞM����vT�Њ�!��A(K��ߒ��:��ٱ��e��w��ӓC-&�:��/�=��3w��i/<]���嘆�[��[u:G���Άgw�4���g��԰$��P�����Ū^�wQ}����K�ԇ>�Zݻ\��0������(�5%co��7�c�����$�C�(p��RA�$V��
���Z�b2�n����N�x��`@��y��N��p|Q~800�F�Fj�Yzw�cM��Yg�Yv�T���!O�3�2x�nb@Gm)S�:�ώ�@_ ��_v}i&��EѺ3I�h�\$�&F`@2?�ϣ%lWZ�kh��f;D�@���RɴLy֟�V��/�����nW*�$��L��/5\p�}2N����L~��Mmf)EB���H0a��o�n���%`���<cwk�T�'Nݍ3ҽN�g�:5�,�K|��~����5���� G���B[��e���D��=+�@���X0&r]��\h�DHF8hm�|O�Ü�aB[��I��C���ܶȹ	�[�;�;Fr�GD�ճH�]
u����M��N�gC��L��RC�=��X�̉Ξ�]� ,S�r���72tW��� 2{@�9�:B���>e_G K��%�n2[�{L]bb�9+UC���܇xr)Cp��ᐘ��zt.`Ո�t�8�B�|�1!��>�	��s�c������Avn����Q�(i�3%���Y¿���p�6�b��)���N���2H.�LK� �`u�\��I������n�eҖ�"��l�lALi	��"{O�'��fR�gK�=d�%���$� +d-`�n�&*7��D�oq�BRx,*�lkD����;͆X��JY�Fn�.��-eOwR��"��3�LT��=���:���,P-��n,��U�| QdH=f��T>zT`��ǌH%����� d��66�V���I2{���+��y����˳�цrG�$b&�v�F/��Z����������������f�M��1��|�����X�rrZ�ɜrV��{;Vl:y'̠t@��E&�E	*��lŀ��8�5��C��l��b��d8x�l�t!`�^^�j����^����������o�����>]�N>���vWW�U=xtU~�������{��V��O뫿��O�;�-�>S���,��wY��W~�����:^ܭ����w�MЈ���F@�l����FFf(2p��L��Y�̈� �9�zQn46�P�jI�1��я2]��%�l*f@:Sm�\ ���8����;���`v��<Z<�ԁ0`v�+'+�[6b+�wPH�7�yj_�5����
n28.Vo�!3]-G�&�M������g2v��y��5E���g�%ǎӬ'w׵ć�5�}.<31Hv�.Sd���Ji��������T|��rn�br�ŉ *A*$��mݽ5���������\����z������B�f�^��:�^����DJ��|x��q6u��ԽG�������G^�W/����_nj�&G�y-�Tj ʱѡ֙�l��eg�7��1yc��N$���#ҵ1�4�q�$TB��K6;���:��x�ʦ$fN3��I�"�(���A]�:�H�]��{$�#�@�w�K��<�&�F'f�8��vi�A�n{��:��ˆ�z6<��Q`����J
���G�dۑ( t0�9�*�T*����[�����|�V��2�C�ւ�HWX근����z:���Ĕ י��5�����6a�u�0<�5�,���-�Ҍ���|�%�$���Ȕ�aiY�0��������ɦ��h���ҸÝod��x�]Oa/ES2h`K�:���+��z�H��N�@$���l�=.I�R�שg>��^AS��?���|�ɎDm�"�A�5!#�p�,T�����_��
�[i��RcP����{M�Ѯo�bX��+p��&>f��t�^��f�<~c�i�~�1j�Չ��?���Y��uQ����,�8�{��9W7T4|^��� 2ɕ�
��K�2��k�C�D�h~$�''��k+e�}'t�r�!'�ށj䞱�K�sRӪ�Y2���8�=����+4�4��g��&���غ���{���l�_1�8Hu�M��3��4�L��{'>a,IoA�0��@�Π!�i{_Ѿ�H"��� �4��-f3-o'���v��RS�H�֍�R̪���X�W�������M�fH:,����c&Ї�,� 5��H��:R5wD�K�B8�S\ R,�����v��2����`�vd˭�4#n؁׉ڟ�Dm0D/�L2nYzԜ.�k����������������~j��_��'�����EgLL�^�mו����{KP��?��`�qt�ݭ7�a)*�7$� �sHBmhġ�&��dZ���Y-t��H����jUg�C=}>���
�De������Wۺ�Z�]8	Z!3��S�g� 3?=�����䛏��źNo?S����$_�q����G� �vh����0��qd��G�Z2Iqt�B�A*�˸�	�t|ݬ����:3�d�K������4i�Z�7`J��-��<��'��7��	���3C#���5oR09�����ЛH�j`j'߲y�)1N����v��8;Í+"��0�Zsl� }$�h&V���hf��p&1З�͐�!s$Y���P������f�M=}>�g�:�矾So{��z�٧�٧���35@��r�CM�Fܭ�M/��L�f��8��j[�����bIP����������k��r��?蔌��膨�,��$~df�p��1G��*ӭ_�5�\�`�9d��,!M��r���7)��~镪w@��e���4���@�s���"#��Z��Q��K����Ȍ$>:�d���w��!��)	t߮��ƚў��e�y��NH���<��O�k�HƱ�1M���[�A�7>c��� ����Glƥ{����p ������͵t����t9Ȧ컻�$@>�{L�5��k<k2�
���R�&�l�ލo�4IAJ>����f����ڳz-��1�1��q�d��\RW��9�B�O>gܲ����3]W��"���.z�ʴ<��T�̞Y4t����8���y�W���g�95_��O� SO��~n�X��/mn-�
w޶b�כ��Z� mg"3�W{��'�̓�.^�fBW<�kSr�^�wg�	IZ�Iy��z��ֻ wr���ei��E>��<��??}~���4���l^��ٰ�|�c�гs7m퀁U� 6[)�k��ؖIZ����
E�݀���m[�[� � � �Ձ,p�/g(
�?c:�W�7�����̡��)C<wٯ��(]���	R?�g�O��Z��2YB� �+ظ��`�@�2��[�Q$��&f<w>S*��jN�{�w+ީ�L�Pe@�z��3rj��R�iMmFq�]��:���N��Q���:�=vL���a��x(��t$)P���ſ>3]*,�� ��� ��1�~"U�^f�����&3�&����i���2P{yo���O��>�N�@�5�Z�H�ߔ�?">�|Yv'����
qm5r������͍�'�Q�O��ս�j�����g��-��m��׵@���~��������RO*ӏ�+�{~�}�;�^���v���L��R^�܄ ��p�16�V��2����c[J����0woϲ�!��Ҭ8�z�f=��a���ȣ��v�k�h�P�8%��Qfeم+����b!�܅��g���N�yu|0����"���2��̲s�x�@s�c�IYE��1�����aD��4����G�@^����::�bL,Wܨ:k��l��� +lA���bE�4x���	��P���z�CY��t	T���ʁQ�7GKq����@ìu:�A�e�s_s<���F.�x�����3;&v�˞=�̛�,)��*�ъ�`g4dT��3�d�)4�����T��uz���)$��z��z�|�9�OA�{:��|Zg�YMO&$�Ǚ��M� d ���m]]m����z��uݿ\�돯��զ.wu�9����!u�T���&Ȗ��k79aj�(M8���"����z&R�߬dW^5YY�0f�"�d�S����_��]�T{��v�tکul�V�4��}fs�Q	xd��Z��3D_�|(�iI��t���mY����<J��tSNka�`C�� �Q�@�+Pa��"���i� /��F�#$�*�Y;��i�'����d�
l�$
#p�?�����;>�����L
�yD#�lO�(�F1� 	b���;��s��m�bY���(�O��IM���ZN�����Ib���>Z#J��_O�����ٝ�6`J��3�_&Ď�h��{E|pB�xL�4K-����� 1dM�grl�I?-��,�B��f? 5�@�7��yM�-ۯz>�W(��#���c�`���y��(��.>ʰ�A�G�YNi�p#+���`̎�Y�g��SF���ʲ��I�?	j�lM#i��""0BD�H�(K�ۛ�$��ubWg�f���o��7��׷���A���T��H�u�9��(Yb�D�t�d5?��.Ky�6�+�\7b^�-}�i���-�����}�7��6����^�|�N    IDAT!��b�Q{��9�>*�`�&K[�zz6���S�B��o�`0���g#��>� z�M�K̘�fxDP�.KC(�TxM"�:�e�bG}��`�ecɼ�B
	��5bqfs��FP
5�m�`�B���P5�Ϥ��*�A�߁���fԭ�Q�@�#{=�����1q׿��W�i�7P��Z/	���l܁$�`���|�l.�cb1gJ�u,��HN�e�T1YB�g�1��!f+��$��H�_�ͮ����_�&�)z�)}�s�8���%�����z�7}u����fL��꺍v����1��/ݯ���eW���Ÿ^˙,I�tQf���-\�)��S��O��
V�&����u���k���=3�S:0d4���1dE�j�]�d��I���2��<F�KnM( ����'^���.�z�d4[�`�.�;�J��O��Oc�J�)es {�"��^�G�gI��h�u�&H��I�Bƣ���Ә����<qCb�]�ӛ�A�f��0"��[0���c2/D�ڠ��r��[ݍ�~� ��d��=*�,6�"7LJ��@�1�64!$8s����ƣL���82�jEÏ{J��
ɪ2Xh2��|�R�B��3� m��q��.�"#�z6���q�)e����VT�Ύ��ټ泓:]�LQ{
�5km�@��@��q��嶮W�� 0]՛�z����f_�H�N *>fƑ'�D���	�Q	�` b��g�$��Pk��m#.��[,��y#r7�l�D3YҤ�ir���e1��� 8ٮVg�q���hy����a�Y�!���r�qQ8���#�L���04
p�ob��"�~Y��l��Dޔ|&s�,�����MX}L�g*㵍���Q`b�,l��rv�N����e�>�!F���#�oiձ-"�6 ���5�"&sn�`��6�e�h�r��-���X�m)���e]�������
npM ��+����f}"-e���-�L�C�[�'n�bd�������=�7;2[u��`�H�2H���u��Fp�Mڵ�NS�{lzo�dV��#`J�tlb�!!�]uC?�JC��_>H6G��9�������ZP&?��Z~;@Ft�n�'EcFGYe�U��Z��ϳ��j�o���:��s}\���e�8Q��Rn�Aг��_�h�Y2�|V.�jcT�M)�>܇�?�Q��ƭ8�2��a��P�]�՚J�$�O�"S�O"=���κ?�����j��ӕE�:dԭ�4����L!�j+�������Q�n� ����u�v�ygH#�:���w8.J.�� � �U���e��T(c�x|w�1� )3����kZ�R��w-Q������h����]�k��@���$�0)��~��$��ݙ�	5����o[a�#��D,�x�@L�jWp����K(c��왈[�����ܵ�G��!��f�� ѧ�4��t7���-�lX9�$��O S$@dsL$�l�v��/čՁl%�8*�*<�&�|��qm�#����s|o{��&0^�mm���8�j��W��ƞ1�#�)jL_|����O��~�c������A�9�qӴ;��Rm`�����5��5[���66�r��Ǐ/<6ą�P���� ��Xf֚z>���9�bG��TFF���p+s��������B�� ��9%V̼�:�ݖNJƄ�)t�#�l(��������Cp�-���~$$��~(���_ǧ�V�	����G�V���?r����	�s8شU��F;τƓ�|0���Pk0��Qɚ6��ϭ�^�V����}��ʮ�Zۛ���uNF&���`��%n�
��l���^]�OdVu���`M27�q�Uc�*� 0�s�\n��7��֮NO�jy�d�h���yv��6@����`� ��T�]&���\��r���z���d�Gǵ�5:�Puߖ�ts*��04��u�l�1�5���)G�� �ǫ�`6y��EY��Z?�XCE�g�7P�=�G*(��2�C�s�/�C�O<�1#$�H� &K]S���{Ӟ��t�l�@�j�Q�ps�F���Z�E��3� =ɹTD�c�45}z�����$~Ί�CNi@�{s�;�L����7�k˨*�x��S�g��P�-f_�A�@P�;�=J�G"c���y�n!���7����"�?j�h�}�
�7dM8ʮ�Y��1���������j���h����  e�W��T��NF@�[��oR�N�5�����f�:��sM��=�ee�>��
ػ���`�ǯ!���إ+<�+M��n���d[h��=�k�e��	`,�m��#;^>�qcc��ι�p_�!�탆���}�o:���N�Rـ���7f|ǐF:?m��;��;�G�!ζ7���x=G�x1d_;A�X!׵��yS1hDk�L.f?R��}�{Y���W��c<�P�^z��7@�l�ٳ��6H1��Mֲ�Q�i^;:��K�¶.�v��;�l[�k�d"��]+������P:q��'��mF�9�|��&���p���;��aoD%Y��&R}�����A��?����ׁ�i{$�|�wW,� �&G�ʓ��	�ҮB�Y~'�F�I�GCWz��� ���j�{��'��
1�	BR���t�7�O>��C��]�8�'t��j���Ό7�hВg�s*��X�to��P���. TD��l�bE�����I߇\ݖ@������خkg)�b�f��o�����Ԛ����7��G�o������W?�j]բ�;uF`du�-������jH(�e�beLa��p��o�����c��
^]^��KS�6���'��y�:t��P��\�{�@��)�����8wn h��Y|�˙���Qh9R���9krx�?�)�T����2� :�^E�̍���o���9Y���$]#��+���a���;fT� z����q�ߌ����F�V���fӓ�(E*5�d���aX���� ���i����E���l�7�|�6����� |�f�Y��,��������s�3�co$�p�1�
H�3�J�K'�e�\�';���Y���d�iRw����y�����#p�&��{/�T�[|c,f�6�Zn���������	��{:�grR�m(�h���H�! !߉��މ�;��	n���\�v����z�r?�::n[wR�-�����+�8�U2�c���;�|�3cuM������~� 3B��v.u�=wO�r�fq/�.���`�I��@���ȸ:������qH�$�k���Өc`�e�|�,s��B�bvc7G�c����_ 
:8��˞�i�j	T�(#h�u�~�;���z�F{0v�	,�ULb�nw�4M���@���+K͵i�`��t�v�,�*$�U �C����N>S۷��k;P��?)f�}����9� ɀ���z;��"ݡ���t�~1��8KքF@�2ז_��y�Ė�I�K#��>�t7�[�g���,�8�+waw
IҚˆkF�3�	��W��,5G/��y�$���W����'$�ɧ��o�n�l_�l�wJ#l�١�gC�(�X#���cWZ�(�\����|uG.e`@�M`��y׽ëb!�]����g���h�X���q��a�mg=�Ǫ� ��_����C�����M3͑�~������a�-��fC�k��i{(�
E�xQ��G���40� Q�Mu=�#P������IW�Dzo4p�6C?g�Z��S�$=VR��g:��Pߐ4�Qs8��$M
���$�p���%��G5�U�&����XE��!I�]m�Xſ%��|ց&v�$Q���q1"b��������b���9���8�\s7����JY@�?�7TS*S�l2��6�T����^]b �3�Lm�b�)'��;�/���)��K���N�@�� 0]]�Ⱜ�����z��~�L���?�Տ����_~�KuY��>���3.S�dJ�S�>7�b���#/.�
2ÙU�6Z�Z��m]_/[S� I�%�\�9��>T�g�U�#5��]V�/�3�^���1������0L�qA��k
��,������7p��Ħ=K*�I�Asl�f7�b���������Y�Ц�Z˂40*~R�Ӷ��*�i�0�g�V��7ƛ��ƹ���G�S����1���k|�:���C���G
^�Q�#-Psp#"@F�]'�J��Q$Z-Y�%9f��=�ӨJ"�ן���s�<��N	�1�'cF��؝�l���N�3n7�ʏX�z�� $�Q�#�����昫�דPS+}H�6�]��W-�2" r[4�cf�ݦwGǵ�GA�:��#KǣrOp �IH,���w�1	 �8iõu�"�u�r�	���ҿ��lt�zF=K���N�����M���p�r:�A���;�߄��	R�Á�v��\��i1�����~�$6�fp{�0��zv3�=RE��x�9Ʊ���BՁ��}�6J����]0M�O=�����b��'�eI7���jUo0�`��'i��]�6ӾWp"�J<2��I����(p��o��7�zF�������2ׯ�F�+�.5�����w����iz��|ٮ)�щ����#�ɸ�t��jd�;�
��C�ήi``$f��rNc��:Ǟ�k�%�/t�!��Y՞�׏4~X{!��C���{���z�Vps�lG�on�5�/�ƭ�4O��ܚ�8�	ٜ�mC6�⻣>�|�gl�����h����H�e�*���d���t�cSQ��K�1��!}�o 2�w���	&Jy�l\�� �MSB�J��{�mhd+��c:6��>��B"��X�1�i�ρ�o�IH	�ɇ����r4k��:k�r�Ap�^���,�.�*�]�+"������7�;�LM��ꥉ7Ս=�7���d�	���g#� �s2mR�@:��Y$�@Zߧ9���c�>��H�c���]��Q� ��\]��DO�X{��'��tB�œ�E�"��s�'Q�X�x���i��h��g�w��� C�}%:��E��|�O��IF�{-J9>_f�U��յvU��|��I֖�r���q�Z����Ds�-cj�#��|x	Rj���fU��U�m��_�3_Q���?Ō������u�{���������֓��`��ZMҔ^d�2����#b��A�� f���{��Z�gfa"=��a񮖄��hL��%6��7���qxJ��[�v�svF�=j���l)�5��V�=7� U��i��<�2q{�I
7�7YF���N�.��$Ӏ�lu���x�`6�;�XX�J���lp�����ӛ�f�҂.f�v�e���G��`��3�j2^-;t5f�*6�A���Ƅ'��')�jl�F�e�=�$���@ꨦS����d��d��I��g\ϩ(��OΘP��a��3�L�e�\O�����P!�AR7꩐��0���F�d�p����u(Ij 	 ���ɬ 3 J��X��Ҫ��E ȸ�qz�TS�@�g��,]U�$��P�� �.>�.�(6n�?tn�]�/L�1���(K5CM���{o��gsc�c�$�&P��ɿF��'�m���#ǫ��ح4]J�(�`�E�5u]	�xN �݉4�9Y}�)��)͌�&#d"�	Xl�*wB3ʩ�Sc�����bʚ���r�A��*>�8A�_k�c�ɵcf�O�sCcd�js�,�0�BpAg�g��(��� �'2����@'R�AC�e��Kׅ@^`qPǴN�����)�����' 	��3P⺏w�sD��dN�(�ݼ>�$'2C<K����:pt3����N����F4Ds�>^���Ho��.�zh�1PQ��K6 ��LI>K����g8䑇�i�F��=�[���{CJ)p6y� ��l)gd�RΤ�Wo��8���΀"�FxV����B�g$�9�l�"R���&7���g���8	�u�?4�S�;)�+i��5E� �R�����Q��rMư]��������V���� �N��!�Z�.�����ۑ��݁��.��V�������s��u��1�Y7gA�D,8X�����g#�<m;���s3��� (f�;��+Q�8K��,jB5Ə"z�Y�o�y�G�1N���'A����\ň�]mX�K������b�����wH�=����4��j(����V弅s�g���#���P<)<�'�̐]H̙dӺu����/*=�aX�
�@ޕ3�]g��Z���mk�ìߨ�\�f��fٳ���}��p]�:ï�Ĕ(~��v�Mē�3	���2�B���]�����:=,�|����O~Y��|k=��Hy�7WU���W?��~�l��ƸfM]<�ntb��4�X|u�L7A;;�E�.���ʸ �cX�bybVU��dKN�������z���k���V�`|_lS��e��͙�	xN�F՚~�����G7�mk:���i���赝��fsF���P��:��g46���^a�(&Ts̰X�.�",O=��<��	�-PN@�X�;�����		M��*˦����Ԥ�X��:�Q�,P�aΎk~2����o����rW���+�f���c�km�dm]����8�4FJ>H�b ��c`���M[��ɔ��E��Ջ4vȂ2Pc�k��d�k��R֊��%%(�(�öfS Ww���j�Yך�٘�2���<=�:����]��T(˄�{�Nw�g�q�3�Z4[�=���2bv����dX@'������f���j�DF�H�ל��II���+�W67��<σ*��>���c�r��e%-��\5՛$�a�n\�$�f����Zۮ�ىr�!�p�d���%uJf�ײWWeJ^<eq�-����,2�� ���=��k�fGf����U�&�I���;z(�l�cV\����ws�X�i������:��B���2bXz�ё�e(X�`i�{��5[}�h�`-d�l����[�����d
-9aG.����2M��*!w����f[֨�DjZe�	�}6�y]]#�-�IG�Ie0k��'#�ĭ��Bꮳ���g���0��:�.��#i�}��A�q�˱���n�e�&5#�k',�����?:�ō���,D�'��t"��Mtu�mrF�Q�X�X4֚�f���(jXi �Un���f5x��Yה1�q�_����4���n�r'|�<*�{�����M��&&��g*���B����3����4*��h��JY5�\�h��{������0��5�j��Ő�n���Zͨ�+>����0�Z#��do�f6롎�}�ύ�&u�5�Ω ��d'tP׉M'�� ���Pq����dJ����V�XҐ,{W1b��S��H�,����WL���&hL�vܿ��E����&��mm�5������)��~�lܦ�r�o��{uV0�@6��N�<��`� �Q��~��_���=�I�7"�tͻ��-k?	�`� �j�����n�֊������gT@��?���W�M4u������S
�@b+�M���tr\�͊���n�֟���5��!���jL����վ������W��nR�!�o�I�8"e�1,�qchu����}�f�y�D��B�+9�,4�i�2�M�.�3�6�|�:���/��|1+������-�q���y-�z��m։>����}��z���ڪY� jfqHw�^������{٢;�֜E�kX�a�����a'�8x�57g���ׯ׸/|Ng�x�.,�)���5GU�������8���$���c��L�N3B�Ef���:�զV��Ca?Oق ꘠�N���:LN$ךFo��������`7u��%X ���{3s�͸H4���3{6?���������g}�[�3���z��-�|��ź~�W�?��z����r��m<��fEG���j��j�'?g�}��j��p���k�l�bP#u�|�������z\+��X'����|t�b�'rP�=O�l>��g��I�~���jW�喲y��xf���4=�lb_�sȥ�]3i�  3IDATs4�@L�F'Mg�:F7�颮��z�������#b���:rwD�c_Wݺ}nc����-h���T��ǎ���x{�jLc���p�� H�ٜ�Ζ}2ۗ`�y��K&�5�n��l-?��٨����5T#���e���Vd���Z���A��0��f���t�n� ��L;��&lf�[ o��5`��nI�D]�d8�0s��90��pˀ��r:�y�٥��q��YN��o?-u�:���W����7��{�.���%�73�����*+a��q���E��2�	�Z4�wqF�B�ב���`�l��LA���L�'s� ά]�s�oi��@�j쓅��@ƣ�\d�������RW�I��w-��L$��f����2�� ����.�8P[W��gvӤM�=�%�q"#މ+W�q�R�M|�lJ2n�7�_��y
,�yo'S�օ��O��]z�7�b&T�z���(�}d�.ֈ���g]�3c8�<�����`�����J?�Fr�Y�)��a?5K����ƙ�{� ��}�$�3a��zn�Ɍ�3V
� p�NYb���A���`{u�Ň�g �zd86�U8�ޚ�$��KpK ��f��M��Fs�������`h���!�8�!=e�P,y�/s��a3_�U��!��45�y��r)��	�ViJ@��H-zp���:��u��,�F�x��h�L�Cۯ��(v�����_�S����&��Š]�쪷���#XO��!k�N��ȧ=6Re>R|)����tI�l���R��:So|��7}K�Ch]�YB������H���2�_[�v%����JFD�8�#��"�U�ػ���J�i�"�����P�sz`�>h�����0��fo�5�]֝�����/���T�>��u|�>�K}�q}��{�`�a�Z�k�q*� H2������l,���S�񢍇��:@~�@%ƿ�ߧ�dv���~�q��9�|� ���b����e��K��H䇔�DS��ty��ޞ�L<�j���S�09U_�Y\�` 4Y�e'g�s�Z7�+F�q�5��`�'��J���V�� T�4ű���vg�0x��,�ǘ���46^4��U�~[O�̑{���/I�hi�J��9�uգ�u=xtY+d=��dX����f.�P� ��W�h��xZu
Pz6�g��sO���U�s�Ѝ\5;��7/�^y}Y�أdy5y~2�[󅤱Ƞ[�@�����k��r����I��x�C�oY���Y�����5-&9Ђ�����^n�7ެ����G�ܠx�����3< ԇ�6����z����'?�JmV�� �� �޹��;������z�[u������yMg�u|rB�<�/��<��ރ�z���������誖�]]�D"��>����Z�W��J9���x�XW�Cg<��g�~���9e'�dЮ�W�����!�Xe@�Uw8�Yo�3oP��r]��Jr23
C�Nݶ�j��`8q�;V�SH�I�E޽?�|qZ����t2�c�w��#[���I��%�;h�K�'`X;7�I�&����$"q"p�0p>��ݻ��� ����`V�f[�.���j��=:��X�V�u$��O�]��`dL�5�=��*Ж�e���>�c�Kx_J{(������ґZ#���=�<�:��8��[��<���J�2��`�rA�e���:�?���R��ά��~���_��`E��y�ZnA�N�X��/�y��&I�=��(dH�juE����ty�?�|�oQc���\k��d��3e�?�<o*5,�R`�g��M�4���	�0J*ͥ$PA&���!K�1!̘�vK*b��p%O���+�t�G�WXC�u��0�rʝ���r���������Ե��ö��K��&L]�=ȃ����FP���A7	n��4�b�9�����A�fn��X�=׊��GuK���IU˝��Sj�>���F~)���� �;���X� z�ʠ�L2b9?�؉vF�٧#?�4��AY�V��P���D�H�-i0�R�ZX�$��G����6l�B��u��Ȟ5�dʘ�p	�����P	�TRi�.����wi�I�Z�Mp%	��<��&�����uD�fԃ�yI8�lr�kH31*�,!O��i,���d�Y�{k�~<��l~�\�7g�wY3	l�����#A�ۓ�@��Fu7�����org��_ZM�U/L�$�7����b�Ԉ�����Ü��W��EB/V��}��;2�π�k�Zk�#���z2�qY��P�W(+.%{�Y�Q�E!�̦��\y}�����T�ͺߌ�LiN�C�^G�+e*
�0�gK)�|]��q��w~~����z�S(�Ke$�b�ܷ�kw� @^��!�q�}ı�<�ě럇}���( �s��\d�g����u����7��5���Q�x�l�K��u�M o�l�:����������6��?�A�ss-�E�/�Y��mXS��g�������t�	�ɫcKd��\oc�����$ul��6���C�W����PcL��Y����؏�|/�Ĥj>�:�V�ZT-N�w$碤b�b���B���&�!������̤E�����1��n�<w��ͺ� �<aO�.VU���Z��YJ���Q�A���d�k���x������jśCp�t~6���iݹ5���I���ܙ���[�y�|����zS��bW��Wu��0�}��4I�Ԓ�d܎5F�-�Mr�#�����cDԝ��u�@�?���j�>��G���\#�-�6�.7<�Y�(�����y~�:㑆rRQ�-�{A >[,tH%p��������G���e].W��"D�y:�ԝ۷���Z�k���,f�S�y	� @����J~��׭�Sf�A<�7P6��@;@�f'�Fi]/�X�٢�i�:_��O�����L-� �Y>�{�՛/H=�ZփK��Pݡ (l&@�)'�줍�3�R'u��q/�.���X��f_�/�u}�������F:�GƦu��l>�Qv��..�uq���r����TJ��G��T_l��x�P���t���$��$N5��l��}j�����Z��yN���/���=���_hR�:��.W��^o��z]�Wk����\�(����0Y0��?�ծ�Py젮Ac3������L�Z����M�<�g�lN�.���Ͷ#H��j�b?��<���%�*agt�������uvv:��8@�����ř�����z���&i���w���6m�P�AU�W�z�誶(���Ԏ��t��a� 2gsDu�!�$;��y6���85~Ü�l��9���ͩ�`�_ �5P��2#�FB����Hb��k�3�ײa�r��Eay�%� �����	���M�0J����y�4Z����)CݫeWF�����8 d%��vS�j��n���=g0��V�:I����2���8�Ԑ&�S$<�!�I�
9�DI��WR��w+<�g�AӴL�	6������샜��m�6�&p���R�����Y,��ZC4�̗n]�Ue�E"01�� ?x�{=/�L��l�M'c��W�S�9�kJ�h�P�ڌe:}ίa*�K��c�Q\��
���0�Lm�����-R.���#�VJC%'��
��y|C��+y�c�0D��lYB�qn$B��j
��ǒ~v@�_��%�uʜ^���♻9ߙ+ż�Z��VB4d����Y��="f�4A�*?����J��L�6J��DMF��p���ҿ��d���Ѫζ��[����G��w���U��Y�'?Z��)��Tn�@�eT� N�{r�Q��h0<���_�щQ�4��1�)�ϫt��K��~!f8%��}PJj����Hg�X�>�⒅���=h,|����%�ނ�$�v��P�zK�tp���(wʕ)𑳡�a�qh��-���sK����!X�Dz��Ca۔��I㿉��A�a"����E�f� ��o�)#��}��P0����b����|uv$`zzR5;:��=�Ԍ� -3��@kق���TCo	�����d�z��a]�ƣ�o���0����=E��k�"��{kk�C,@
`���T���c?l����Hrt�X�$9��%W#�v��������ve��@+`�O�An��j_�Ì�`���0X��t 94��d���!C��{�k!k�&�Zc�-}W�>���d�0*6ШM�Fp�u��  �U�}��V��I�b֟0�>�x=H�$ H
X���_̥��ןJ*��������l`���������9�������t���Ԛ�,� #��jf
g��,C&_u6�uf�ˆ}q�PC\_���@�$�L.�;&�Lx�jU]]��+�[�eF"I)��]T3�!cy-�Ꭽ��d��P�$C�cM�Jq��<���Ҿ�n� �"v{��5I�;��{'5O��)�]�UW���p=��$�%5�}&��2���j��5<]7��l�)�KS�
 D&U�M�X,���Ԋ()���1V�������m}.���O߽CB$��Q��պ�x�a]^���jUW��=�^,%S�7"�/��N�2C6� �OvP�iH��ڽ���Z����	3�q��\��P�X2��X��f$�ѧ�[CJ���\��Z�/�G��* T�V�K��n;`��D��׉����"a��o���c�n��5Ȋ7�:���DP��?zX�߫��=iܛ�eV6�SO�-WB-6b�4�L�I�4B�?:'�v���8�Ź��N{��`j�>UN�gP�g�5��2�ͽ`�(��~���8;��z�R<��N���+�*�C��s��,��r�,�Veg�b�l(=�2�RL���RQ�Fd��)Ԓ�e�[3ρK�U��IMz�8¡��#�@��i�=� �?��)`�M����1q��IYaTx[0�T\�1I����(*١dm�� :����D	�˙��k���![��%�0$����9�Y�6�K�ɘ�?�v	=C�:�����м4��	����>	L1Mb~����W�۾����w�H2�mCӓ����vTn#    IEND�B`�PK   �c�W@��-p:  �C  /   images/f73b1f81-ca5e-4eef-b776-593c08c8c802.jpg�wTS]�/�i�ҤW�RU@DDD��J�*MZTP�4�����" E""]z�t�M@z/��B���S������sθg�Ζ1��Z���k�����LǴ�4� ***�����j�?����������?t��(##�Q&f�cL̬�Ǹ���sprr2�p�pq�qpr(��eh����`b`��_~(_���7*E*!��������@ �������PQ�>�?|�(���@MECCMKs�5����tl'eT�ܥr�8�$:����:N����GO������?u�����._�������u�����춹���v���^�>�~���B���x�:.>!�M҇�􌏙�����KJ��+*����[�������������_X\Z�mlnm������ �?�����EMKKCK�����`+-�I�Cl*�w�م�?9�q-:���!��ޣ��\"�Dq�~!�����_���50�P�ɣa��>��3;���'r�1bi�(�̃h���-�Y)P��=)=zUB~]SMڕ�X�a�)��2��7Z(��zY��x�%�ba_�l�vy"�n��}'��
�m2�/��F~�v�����s�ZHޫ��Q�ȆoA���N�Z��
(��M�Qթd-��+���O;������X�e*����O7"�Z�nL}#+ڑ�ȱ�u�)W�*�!nF<��c ��Z!
У�+ s����E^,��U�o\�,t&�_������K&�:o����@�D�8>���7�����6���}���'&礍`�鼭-ej���X�����Mmx��}�ӵ�>�;�ظ��9Ȑ��|����й�/�vg,���q^@���ț��z�h[��7=�fO�)�/�3�j\����-q+�S<���71�8�r:T;��7�t����()2_�K�7�0O�����^+Uϐ�s�)�0� Z��LQ{��\���J��&�\9����W�6� �(�}��u<�ߤ\�/[S��X҃C?��C��]�b�\��of����_R�)|3��������6���#�O����H.�)�C
�����H���R���~�������Y�m`	JC>��3T�iH�p"A-z�OTj>3ep9+�2�*rd�m��@���D�^�3�� ��ie!���GL=��f�'G��^5NiB��T��v��Hknl^Ty�������4@��x4=���G<�H��P�L�)�d&Z�C���?����\ls؍�,g�o8�� ��8;�D7�yt\ �1�7qJ��S�q�JEWįdZ���}�'�eFOE ��%L+�4\�W��h-�~.��*M��H�}9�|�NTvWsN�͂	���q����P���XII��Mc	_nw�
�YN���������;�X����c�/Ua�_���N3dV��3�]T���p��׃�s�,�
��͝��ZN�Fx#�~鍞^m�~/!�5qSö;Eg+�j랝nT��%��  ��py�Y���y�M��������A�xы1�i)J�d��p����8l�fa��������6��j��\+�=pN����HhL�ZW���]ՌJ��`��@�Z�M��1�{�i�N�w�C-QF��v���^�>��T�s���A]�X[�E_�X��l �\�-�ݙ,H�FaSj�3��W�NJ5�ut�1_}�2)�^ak�n-:�	㮆Lw8������{��
c�U�
GN�2���<b14�4h.Z��"]_��7�stT���5���顎����)-g���\Í׊�#�q�M������N���V���_�r�����[0�l��f��gV�y$���f^|ŵA�҂$=�8��A|��I��)��!2W���:���)�%y3��P�0�o>/w����ns��ĳLO�}����.�n)W2E�N|R�:rb��>|�[] ��������.
p�MV��B���\N)���d=���6F�T{֩CwiM�H��5ͯ�� N<��2:�%��+��d�K�W�E���Bi\4����&w��&u����%�}�	
�8��Nk�d�s�f�������֯� ����O�雯���=�e��x,���
l����k����Z[z�"�O1E�e\em�=�Ƣ�i豤�Ѿz,Gs���z9ieT�I�*�����e��E�vf�����[�U�����V4����ng�\��{����g��~�v4�.�a��4�fe�����%�9��K���	l�Hq���Ҋr��;-��e�	C��؝�A"��B�g�r���QdF���}\�-��%���oP-{Raް:ѐ�R9�X���;�5�(��V�^!ym��y;M����Ժ8]�+r/k��E�!��}K�.��3k�P��V�Ε$1�7z~(��O|]�z#����y����@�5+[:o�'��/�{Q�pg�i�ٴ��|�͝
�g�c=w�Fi{7�����ڜ6m,��/�]?����ԥ��lΘ��:� �E���ɯ��Q�yYѻQS�m^0_�W+�.�f������a��fY����!�x����P�Bro�-�>�B���3�c'lR�:\��ՃEqL�fK�?�s��;�-7K+��S��mf7~��$eU��uQ��=x�����f2Y��Y�q���v�0[:�_�.u{�᫓�Bً�C�$����|�Qߧ�e�A�g�!I���-������k&_�>�̥����4��U3=�6�Hڏ�#E�gi�e$[�U�"�I�=�K��Ԁ�!6�WT��9H��|,vPǩ�j�(��e�ba�Y��V1�?�3�B�l癜�W'��X������\\{���$m}��#��R�)+���KN6���[M������D���&o���1�s[�~z`��.�Ȯ�XDF�y�3rn���%�����L�=�|��T��X�Y��D���>�[�o�]�G��t
�o�#W"��DӽD��
��"f�v��7���+)�H��ܷ]��ch�?��?{7���ߖ�ӎi����N:>m2V���?��αo��a�дS�j=ˇs�2_�qf���gL�Й��e��SOE�"���r]����bE9����}���R�SAc�2��gϚ}�i���a�*P�p�����&�,���3+4Y�N�$�|;Y��3�!����׭���])B:<�3����8��p�5�/N�����-���[yɐ)����/��z�*+n��uuz ���+� �UUQ�Cz�5���'��g�w�J��&2�̾��ѝ q��J�>v�&	��$�>���-�LMœ?��L�&�7�?*r)|m�[?Fnz�_�M�+�>)�[����7�:�����h�Y57y����%��2{���;9{9�+y�3^и;3�V����{QӇ.�Rȟ+� QL�|�mN��:�%E��Xyu�ޤ|�0���g~&���C�h����j��JQo��Y:��0�}��8�gܧ���%�b����b�tK��*6�Uo�oY9�:�����)l�'����D]<f2��#���@�kxi=�V�,�Z-�g������K�g�
z���Ja�7�$g�cr`�1��P冎�w��H*yG�?L�w%0`r���Z��H��Ȗ���n��Lu�.�=�4U�^�M�#���M�;o��kpF�+,Կ3+�����+=�l�����f:f���׍�&{�`��|�!/qA}�܂��}��8�itY0���g����l��Xf�#��[P"��^�t(Y���K�FC�m�l�܅�/6���[P�I�l��2�>�G�>}-PP��0��r:���4��O:��5//ݤ�����V��=��+;�|�Ov�g�M؝( ��t#�xi`\�RF���3�����Sg_�+0������pA&��� W�Rғ�tߐl�t�4$��Mj�7*�:o�"���:�1�i���6�I���6d-f�R`9h�
L���>�6k�8�i�*gm-��r��E��Da��0ݮX���7 ՞#*����[��4�޶���}�*!)�^���UO�c�浶�S�����9��p�S��v!e�C�P�×.] 4B^=nt�7�/�oVH����hz�k���
����á�뺎/���'m���҈S''/�	=��q�.��o�<:k��t�� +O�p�x���jWe��}��eM�}�@���U��9���}$s}r��m�,������{D�b�ISs28�>? �۫�W'�Pٖ�b�p��&�O߄:�h�fy=�����y�"��7%%���pX1tu�=�O�d���	�F�����Pm��s�����y���I�`�^�m݈UrM):4����(���O �Po5QR���+�C
��{P�q�0C2U/y�F�v�,a�YҜ�dLA	L����)X��.�˕��C�mIQk�Q9cfcM"7�h��a(�Ȍ���x�Zv
��8��D�������3º��s�o]rq��*/���8�U4]������U�ﰇ�4�X`���=��un�z�f[r���N>;�|v*�nIS�C�b����鈥�(ܕ-���؝���.��d6!�|B�Ӆ���bإ��&�����}��Tϰ����b`�mM��mw	v�0�Ty�z��^\ؔ��u0F|g�l|_�oV�S�܅�0�����WV��'m���xj�����]z�g��y�M(Sġ��c"ggJ�#�G�]'1�Y�s|<ߖ<�,�فlG(|�%6�uć���ĐHy.䬶֔�k��-{ ؈c9	\Ɔ�E-�7Lq~�N�:��i59t�{ȼ����N�����[�1<���*�5�sd�{������n`QZ�S�2���M���3o���ܔ�+z�d8�j��A/���<3άإ�S �G�/9FGrW ����O�w�`�}��%ج�Z��z���z��s���P�N���lu�E����3�5S�*���X�}���)�
�Ķ����X�Zu xJ{K�)&����|_4-I��Y�N�%��װOAC_*z3�L6v˪��I���x�q6��\�>>E{
�G=�B~�U�� ',\S)@w��?��맦�	�=
��Z��"�	�X��W��Lj��酄=u��R�p���f�%�V��u����i8�v.�]Wܹ�~���f��>)E��jtIg����q�1��W�D�{ʙ"�򙊦�;�2�h�K"�`ΔG�Ř
s�ET�$��m����Y��;�:�j�&��x�x=��m���\en���˷�f,�E�]���5�Mf��%�'��:$\�w��5}{�bU�N<���`�}������Z1�M�_�;�oj����Tu�l�	²<Ij^�Z��8���RU��˹W��uf=�y�;/�*0����	�=�(���ym��Ҕ��%��o+�kY$\1�7�Q�F�oMPUK�9/$�n�x������H�������;��{�P	>���ؖ��Ò5Ӑ���T��a�O�����-�{߭~P7t�g�I�~P��[+	�ĉ6g��t�5���]��=0���9_�#��X��T�u�H�g4B`:�kiDq�Oh����w�=�>:G��[�m쩲�X��ݗ�4Q�Ḗi����x[�po	&O�!�|-�zI�v���F�ؠ۱��)�iy̑��ɇ�j�Ԗ�ڨA�.Z6���6����w�t�'ޛUN*h��ؿTzi���[��)�N�óe�S_��w<t�uyZ_�=�����4&r�e�l�!�T���r8�&N;��0��՞0[q%J� �>(�W��2����E�rp_is�^�e'�#�pD1��ޙ_
m(�~q�Ae$�(Ց/���1�z_.�`W�(+���AC�����>&�����hZV0�SQ��4Zw>bR�9�.�������GX�SKJ�zn�Z��-��4%k�B% �u+jU��܎;}�>�D�NVӀ��D(�J���vh�����Q�o#�-�ۃ	���0��rT�d�fڍ��Y��؜�
�>������S7��1��ⴓ���o��z�_�D"mG+U�ey�̭���7i�����զe���3�D��]���������ǌ������/�os<���{��[�!���?b�C�f��W�H�rQ�)�Ẇ?��սXHЧ�E6Q �0����oSAN|�Ӵ�М�K)�]Għ��yf��_4Nl�]j%���+*LՈk*�pUnp`*��X������k<�)�i��dV�bi34y��ɔ�q��ʭ�2�&&�{���/$+j��'+/+Q ��M�
�"FoRY���<cǠ��]30�L�1m�������9�4�N��;�w,���+١;��n�D�B�Q aC9�G��7�q��[���;�u^[��=�K:��=3��M/�0���dH���K��j/��ţpl�`�|����'��Ԓv+�S��±#'+�]N]gjz�ӦV�G�坧�&G�w}��FHlsyI%��>��)��М���fA/a���2咀KkHa������Ԗ7���i�4�N��˔e)@�e�86k�$ҵI^��W������"]�-�k��y�4ȭc��0����=�x�,����y���z�}���U�D��C��b5Q�9���,U{XM��b>L�U͙�j�R:ۜ��3b�=&��Y=��(�|ތ�B�\��	/�w���j�Rs��EU�����Ge[���
���h%c\�7p�|��0����KX;��<�4�۬��3�χ]m�*&�:P �9
0Qgipŋ!X��-|L�_�G����<׶h7��/}�4u�Q���=Ml��t2��9�"����열��m���=��5��Re�ퟴ��� �h�>N�6�(��`�p��-��U�7V��S@�s��\�Ea�"�7,"�������MT��K�Q[,23c;���j�]�K<�AbA_���4v|��)"8s'�V?w�3��㞒��[K,"x�]�*��p�؋ )��$�6�դ�l'¯��V��Nl��f��	M���	ubd�s�M��]��:�6`�'�j�^(�*}M���� Sfj9��j�Iz*t���4�����EM��ĎŃ��+o�ϵ��x�V,;�\�9�=lA�vޅm(��Z9�B���q�2�QX�(z���M�W�N���VA�\�t�e���:>�1�#�RQ�`���)�ar��XI�!Q��fj�f�/�����йbR��Y���F��6:l*�w֋G1����q��F*�d�|P���ޙȞW�J�!x�z�/����[�7�����1�p~��:���OB�uiܱ�ot�4��w��<�|w�:/���bnl"�i�,�6�=��T���JV��Y�ݿ����<̳���L�q�+�����z�V�	��c'�'�����_��;:n~N�I��C�z�/��7�M�o�[w��K�\�<����]?V�:I\����e����Ti;ڷ����"�z���ZK���R�O�Ϡ�q?]1p����7J�"@S������۰�Gz�ɉ�$kwdI퐧���@ߪmwix��2�c�7����ˢ�:gR|7�#&
�O�E��ؖgr�M{̴��?uxW%VT'�q_�p�)vwf�����fm�����L�0{(ޠvD�TW=��(x�G��t���+�2p�]��I����y�r�pFd��7|�$�ٴ[���V$��� UT���ڧ)pO3¾׫U��yw�6љ<�!J�m��d{�Uf������X`L�r�_{}���2^���ޜx�f)9n�8�������qD3�An�ӭ��0e�Oڢ����%�ix=�!��՛��ykzgq��<���h۪h�ai�
3Ŧ��������E��ɓ�0�g�h-�h�)�.�L��N[�a�@���$��{��aӦ<ҥH^|7p�Ő���9��2Ϫ����l��cӐ���j��ƒ���.�s1N��ͳ�����<�sT���e�9��ъ�k|�Ü�"��i��������,_5�C�!�G����:���-"�l:�~����l���W�,YE��!_��7��8�S��E����2�ة���

0�����>w|�g`=�Eԕ��`��˰P�
W��.�z���P��v�4���S��NH2T�0�`�R [���ؘ�$�E��Mz�]��!�66�(�D/�N���~� }��WR��z�̈��
��݉�Z��g�S��>x<r��וP�C�$��5@���Q���
 I�T�eC��46�|�Jz�K� û�@��<�/�;�,�H�1R��D�6�� ވ"�B_�pf�R,n�D�NF�� Ġ���\3��5����,�JP秖�P��_n��M��7:_�_^�]rd�#$��J����R�:����Kt�~Q�՘TZ{�^��I���,J��u�a�࢒[�Q��$���b��A��}{�ZO���۽��Z�����������!`E��GJl�#����uj��]�ѭN1撉W4cg~R�uC9/�]1��L.�1��(���,�e�I3��6vb�i7������Tܬ<�|��y��O����/�+6�Nl��Oy�ӵf=%Y���jĹƺ�~�{}Ηw�Nw�cD�.-Xvn���lM�*R�j���%�*��D�g��6��V����ӻ�-��P	璖�dsMH�.���$X���$n�������ި�k���r�A�z9�2��P�����?C��%�9�F�*���	чE.�[���f�NaQt歹��.�|f�Z������Z1�CMs���V�31�m���:=���S�i�i��bp-"}t�;:��tv�M���ͽI������s���u��=ii�j�P���_�ƹ�eq����^�p	��/(�� ^�����������}.��x@r&��9���H�{�8�+������������y���!���Pma�ұ�0ɒHA���`�:�:?��t�KD���>=���ě5w]�&i鴱�6H	�Fz���'�N'��Z�҄"ʌ�/I�Q�z����\�LE^��GU�9��h�䜮k��!�G�&꫶�C׼,P��ʟ�(N�6���V��lD�d
q+�|�?e�?dk���<f.:]�╏2�	g�A��(R�N���s�+b����`��	6����gf��;-�`k��@���B\��c��%��<E�_�*cJ�󘜜g;�|ч�`ms�Y\�E��+����
c�:���|y_�0˼s�:�1�Ād�M�s����ci��V0�;�Z>a���+����?�ʄ�|�N�Pi�%�����#pY�t�)���c�'�c�D�+(Wb,�e"�$Zm��5�D��/J�j6�j(���#�Nkx�
S�]��Kؠ_�蝹���ז�}s׏,w/���}�?�Ѕ.�i����Ы�J��E5��\��%;-��.�y��~�B�p��r��G݆Vv�vڷHfo26��XaQ�4����H�q���ZLy�Q��o����3S�W��9��V�k��ˮ�F��Iν��W6�{<�#�d�{PC����ʛϼ��&	}��D�h��f��OR�rJ�P�t���L	YDu�g��r�gT�|fQ�"3�̫g�~��s-�c�&U��*�0G�N����7��c3`Y�m�k�Ý
X>&pee�qxǏJu4�=��K�)��si6�	C��5���͓�m��8U�}7ٕgm�+s�v� ;���y��p|b�Ƿ�"A��u,�lCif�%�}�%L���'B��JR�s41�=�9�v���cs�8,��ع�3�Й�<��U�P��X��ә71=Дܔ�$�]��{����ڥ��dw��Rv9�;��3Fi�+�(�[�ƽ=�f�.���\��v�ݷ�7[����[wy���6._���x������X?�]7�p|k�^���W�͏�_;���y��7�m��X�/��,J
V���Q^�*q��E��(f%�n�ek��z>'Ǫ����Q7���\#1��2K*=��!V9���RVA�'ۙ_�L��8�&7��m����J���-0ˡo���p�i�n8�,˪�wOsU8/O;E�7�r�:S�^x.�TS��n�|���ϼ�?mY��]�7��b�����ʅ�7H��N�� ǈ�V�ӰS��r�>��j}m:)b���T�Pt3����(�J���1��������p֬@�t|��ˠ=�����wO�?$)Y�s2r��[�OL��uH��^oe8M��������� Dy��_�s��0�#�:�ȑ�xX3���;|�j'GtU?���j���l�U�݂J��o���H�s�|�3�����Rl��rPk�Y�V��k�\�W7�jYv�����z�����R	�]G��3c殬?����u~0����K��ʉ�m��(,�7q�8bZ�A�x=�=]��a��+�p�ΛEO��|Ie�9�5sM��U>�H����b���� ��;GĖ`5Ȧ�!���=_rK�=]J���
�/� �i���`�R?XT� O\�P�vEݥ W����z���X� B�������.������C�C���X)
��O��]�)�{��YD3R���������V;{���GB�@ʨN#$��]�y���-Է�Q��'5�Y�#0XGjA*�2�Ed@���������zt6W���{\�����)X�A��S���R�T��<�;�D�����"	�U|�(@�s��{�PO�)��QCp;f�L�����@���������G��a�MZ�n	|�'Ԯ��!�}�y�:��s�у�&�U!I�g) ��������(����cݙ)�D���n�NN@�9�����:>:g<��C�5E��>I&K$=,7��?���һ�㷢�N�aٺ_n�ű�5��S��.{u�Ȭ)��r�� ������K�h����%��S�İ2�v+�U���~\��7��(�Ч��t��z>�k�	��}���E��H��#k�A����SD���zQzS����R�^v%�1���ҙUe!��>���҇*�_�g�X~����2�M�i!����������ͤwaS�h��O
�ypb��dR�?5�3}��Y�n��n���ջ�K�K��Ɉ�'ы�)C�4$uS��k�ͪ�����)ڤr��A���0��hP�;�M���A���W�>�y��NQ �yR�s�k�+��N��(@X�w�����kx��k��M��f�����2��S��w�1�'N�a!�yE�rCt?�#��!�iĉD��]�[�],p�"�E��Or�hl���[���1����ux~��z�	<���`C��9
0������%�xP �_@~yν�}�/�?���]�5�<x�ᙡ�l8Cb��o�?]G��'!���K0l������K�N!�K"��@�:����'���_��ϜL?1��2� ��@o�f�=rO=��ɮ+�Q�~4<�~p�F�ه�&�I��9u(@�,�QE&�y@���q݉��Cӓ�Q�1��l��p��
D�	�P���\��`��\c1��!{������*�(@bb�	X���SMȽ��$<�������e��=�&�oszx�
Э�^���D�f�'�K>�:�ЍK��P{_naSd(��E
�sv�m�v�LD�!��<�/���ռ8���~0�;��Ͳ�1�&��eH���!?I�M#�ȳ����4d�'fm�����[\'1��'����p3��Na9P"�� ?!&`VF�j����ki&ɾ�}>�:0�2�6i!W�opnb��dU'a��ċ m�X�޾|�t�9<4�]*�R�O���	�������2�@�Ju /��N�m=�/{����%� :ח<�1�s�k�a~ô(Nv��q�	��u
��n�����L��(�T�$I��w��������S,��R�+��pG½Z;<ȇD�)@� ��1�$�|fKQ���Gl$�Ծi�"�^��k���,�8�9;ղѼ���2�!R�����\��P�b��WxIsL�T���HO��QZv��2w�(!�B�fߊAI�@�'��g����{!j�F:��I�*e5.��n�}J�{�}�CTuޜ�pFZ6VkZ�����D��rIȣk[M6%hO�cy�=��T��s����
��vF���`�+Xl�j�}�f^�9DV�s "���[	<K�?�o�C�/�X�>���V�e���=B�| �J��Gz����]w���E�^5���k�l� �?�(@����� �!lgҿ�*{�z�_WUR_�o}g���\� �|�V����v�?H��K>"7|ѩ��ۋ���c
B|�$]N�"ql�B��j�u�g���#�Ų�IZX��ݜn��L�ަ����M>2|�->��|�!IH���(_H��7�א�f7%�e��f�*�+�-���p�%�'�ۇ*?^x��m���`S0��r$Ȇ`dmצ��UdO�j�������j�>>�0�ˆ�7;�=�3b�>A3�l�w�}�	�!>xK�����FT;���lBz�5�q�UJ(�/�uX&*q{'�P����"�4������˪����@eH��Q�޸ڥ��ڼI�Ft����`O�������������8}���%��u�Ԇ�	��m���1K���+.l%�L�a��_�L��2j~W��2�~����$�K�X겧X|�Xn�����.t��XI���`���*���?ed��\�R�"�f{��t��¯׸��b�Y�ن\�W�A��]�ji��;^�$�A:���������G���u��}H�'�q����m�e��p3(��Z|G{k$�0�d5�`�P[���_�����q��䨛�%��Ǖ(ǃ�s�Ab�ז�"0.C~�Eu�h�����Q<Gla�Q�[P��K��Bf�s%s��4(�#&`�U	X'	��2��j�����f��z0��d�i`S|_�K�E��;�Z1(��K$����s�(�6�S� �`�B�����R`b��{�N�-������Z� �䭽��q�L��[7��0���p��˯���"I�$:i(�$�#a�V"�pqYi*����r��<��Q���)�����o�;��R$hb�u�F ���@��� ���E<|���fG�g:Y��Z�̦dA~����S�r��oW��K��ƈ��qb��~��.a�9�^=�mx0�@~M"��J��):���*��ߘN��门���N�&���*���`g����[���mk��?!��l0�߷!��X4^cەp�������L0��^��7�Uj</ ����=����q�4+�����g�g��rB�����0c��.�yl���p�3��8	��vCX(��	�w�5�!�)��^���g��U;
 ­^�oQ$����ha��qk��C*W(���Gd�����\�CrA>ro����W�7َ� ۆ���V!_$4v%)�D|��"�L�.���������w&��㶚���j?k���h��D�e!B�T�W����(������2�N���G���!���A�>cЋw]����to��ao�f��-�* n�����;��I��h�8���QDw�����U�������?�[�y�a�Gj4��9��[������ދ��.UG��a��}�4��W����/�F�}�G��Ғ���W��|O��"��qy-"W��!W���g�R��-�ių� ��B$)3*�#I�eM�$��F�}l;s`�⭒b	��K���ծ�u3K�c8�ɮ�mݲ���E���:w���*�R�eO^�G��^�/S�~Q�E�݌�`M��㣨dAe�]�i�Ft�k��<{��ؼ���Ǻe�z� #�B��ΜR�5"6�]2?�_�u��=�=
� ��z���N<��@��D��d�)�
�]"x
r�&��Mp̄n�����`��6�8��
��3�+�J6�����a`�z�@F̂����T} �b�0j=���I�x�/2���M�>��7�$b��@Dr��#id��h�.'S��gj>�$�A�\� -��e�]%�b������ ��3�mw�7���1����_�'������@�.����o�R�;t;�Gd��S:��E�X��~z�~�<1�t�����o84��#�7"
�φ�C>���i��� d� �A���e
�c��O�����.#�g���������Y�|�>}�F���;:ԅ�U������s�/���#��� ����Ѥ� NQ����w����@��0A�'�ރD�X���p���$�q�E�9��_xi �3H������9�e��쐡�+.f�(��&쐟�t�Qϋ�.;������:%ƜW�8���|TJ�S�XL�7*�bV*R��9#Ο�T"{EZm�1�LAw����X��k%�6���;�9��� wg�
����!��2�!�8>T���3�UwI������PoO�(������ �h����M����a01�,��� ��n�g:Lu~���
tk'Ǥ>�\�=�T����L�ŮT?��B2�����6�zB���.woO�I|hi��]��t;�n��Oat�7O�C�*�	Q����N3ji�J��T�x|�ԇ'/�%::p��(Sb����ʡ��XvFMT���/q�{�؄�l�aE|۩��.O��O���Y`�U^aLqSW�J<��� ���IlI4�1@>� ������kKMI���~/����ѿ��g�"��=�=�Rcw���B�,zՇl}�*r�%��������PK   y�:X�F?�  �     jsons/user_defined.json��]o�0��ʔkl�����HS�m���j�*�v:Oi�%�����sJ�L!�!�+b����x̖����٪���E���f��v��� ��x�[���.��x�~�ln�ڶ��8Ϛ�����8/����ЫY\��a���0�,PDj�6�-)���7�-�/ەߵ��mC�����ڗ`�nb]������cV�n�kJs^��3B U��8�e첾��0��HN7�͊���{[�.��e"?.]?��B��P�+*����3�8�3�CB���?�6Voo�4�����0����0e��&�l5�M��r*����&��8[Le�q6�ʖ�l�̾z��&)�B��:^j�Ʒ��	��uu���7K�ڸk��2%J������0�\��BWp�r�}!Ȅ(I��D	�I!E	����O�J��Q)a�Ƨ�=%J��}����j�u2�>��=:I�+x�C�?�/R�.$�q�0��{��/@.� \S���o4E�<�ռ�6�\��jc
Q\}���C�(��1�gZ0��"�D���f��x�}��{p<>����;?V�d+�Z��ޝ�|K J1�(o��MY|H���b�99/�)��`x
>�pE|�C�H�������:1�Q\�ٯ@�:{�&�K{�����;�*����iLXU`p\�r����c�;R�	v(�	b�`�!�1��x=v;H��X.�̎Z����Ė��ڞ,^򮭯�PK
   y�:Xp:�  ��                   cirkitFile.jsonPK
   �{&X��N���  L�  /               images/3e5d0cfe-dbb3-4add-86f8-df5e0b35ef62.pngPK
   ��:X��yD  4E  /             ��  images/68f8dc93-d533-48f6-a1fe-8db98063bd4b.jpgPK
   �:X��S�  �  /             Y�  images/a8eccc96-6934-432b-b3c1-5526b5feafa7.jpgPK
   �y&X�,J  /             0 images/d5a492a1-86e6-438c-8279-421a5a29733e.pngPK
   �c�W@��-p:  �C  /             � images/f73b1f81-ca5e-4eef-b776-593c08c8c802.jpgPK
   y�:X�F?�  �               �Z jsons/user_defined.jsonPK      S  �]   